
module AddRoundKey_InversMi
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  statemt_address1,
  statemt_ce1,
  statemt_we1,
  statemt_d1,
  statemt_q1,
  n,
  word_address0,
  word_ce0,
  word_q0,
  word_address1,
  word_ce1,
  word_q1
);

  parameter ap_ST_fsm_state1 = 14'd1;
  parameter ap_ST_fsm_state2 = 14'd2;
  parameter ap_ST_fsm_state3 = 14'd4;
  parameter ap_ST_fsm_state4 = 14'd8;
  parameter ap_ST_fsm_state5 = 14'd16;
  parameter ap_ST_fsm_state6 = 14'd32;
  parameter ap_ST_fsm_state7 = 14'd64;
  parameter ap_ST_fsm_state8 = 14'd128;
  parameter ap_ST_fsm_state9 = 14'd256;
  parameter ap_ST_fsm_state10 = 14'd512;
  parameter ap_ST_fsm_state11 = 14'd1024;
  parameter ap_ST_fsm_state12 = 14'd2048;
  parameter ap_ST_fsm_state13 = 14'd4096;
  parameter ap_ST_fsm_state14 = 14'd8192;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] statemt_address1;
  output statemt_ce1;
  output statemt_we1;
  output [31:0] statemt_d1;
  input [31:0] statemt_q1;
  input [3:0] n;
  output [8:0] word_address0;
  output word_ce0;
  input [31:0] word_q0;
  output [8:0] word_address1;
  output word_ce1;
  input [31:0] word_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  reg [8:0] word_address0;
  reg word_ce0;
  reg [8:0] word_address1;
  reg word_ce1;
  reg [13:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  wire [31:0] grp_fu_320_p2;
  reg [31:0] reg_352;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state4;
  wire [31:0] grp_fu_326_p2;
  reg [31:0] reg_357;
  wire [5:0] shl_ln511_1_fu_362_p3;
  reg [5:0] shl_ln511_1_reg_1261;
  wire [2:0] j_fu_380_p2;
  reg [2:0] j_reg_1269;
  wire ap_CS_fsm_state2;
  wire [5:0] add_ln511_fu_386_p2;
  reg [5:0] add_ln511_reg_1274;
  wire [0:0] icmp_ln508_fu_374_p2;
  wire [3:0] shl_ln_fu_415_p3;
  reg [3:0] shl_ln_reg_1289;
  reg [4:0] statemt_addr_reg_1295;
  reg [4:0] statemt_addr_16_reg_1300;
  reg [4:0] statemt_addr_17_reg_1315;
  reg [4:0] statemt_addr_18_reg_1320;
  wire [2:0] j_1_fu_490_p2;
  reg [2:0] j_1_reg_1328;
  wire ap_CS_fsm_state6;
  wire [1:0] trunc_ln521_fu_496_p1;
  reg [1:0] trunc_ln521_reg_1333;
  wire [0:0] icmp_ln516_fu_484_p2;
  wire [3:0] shl_ln1_fu_500_p3;
  reg [3:0] shl_ln1_reg_1340;
  wire [2:0] i_3_fu_518_p2;
  reg [2:0] i_3_reg_1348;
  wire ap_CS_fsm_state7;
  wire [63:0] zext_ln444_fu_529_p1;
  reg [63:0] zext_ln444_reg_1353;
  wire [0:0] icmp_ln517_fu_512_p2;
  wire [1:0] trunc_ln457_fu_534_p1;
  reg [1:0] trunc_ln457_reg_1363;
  wire [0:0] icmp_ln445_fu_564_p2;
  reg [0:0] icmp_ln445_reg_1374;
  wire ap_CS_fsm_state8;
  wire [29:0] trunc_ln446_fu_570_p1;
  reg [29:0] trunc_ln446_reg_1379;
  wire [30:0] trunc_ln447_fu_574_p1;
  reg [30:0] trunc_ln447_reg_1384;
  reg [31:0] statemt_load_33_reg_1390;
  wire [30:0] select_ln458_fu_622_p3;
  reg [30:0] select_ln458_reg_1396;
  reg [23:0] tmp_2_reg_1401;
  reg [31:0] statemt_load_34_reg_1416;
  wire ap_CS_fsm_state9;
  wire [30:0] xor_ln477_fu_925_p2;
  reg [30:0] xor_ln477_reg_1421;
  reg [23:0] tmp_7_reg_1427;
  reg [31:0] statemt_load_35_reg_1432;
  wire [30:0] select_ln487_fu_985_p3;
  reg [30:0] select_ln487_reg_1437;
  reg [23:0] tmp_13_reg_1443;
  wire [31:0] xor_ln524_3_fu_1003_p2;
  reg [31:0] xor_ln524_3_reg_1448;
  wire [31:0] xor_ln524_fu_1195_p2;
  reg [31:0] xor_ln524_reg_1453;
  wire ap_CS_fsm_state10;
  wire [2:0] i_fu_1207_p2;
  reg [2:0] i_reg_1461;
  wire ap_CS_fsm_state12;
  wire [3:0] shl_ln2_fu_1217_p3;
  reg [3:0] shl_ln2_reg_1466;
  wire [0:0] icmp_ln527_fu_1201_p2;
  wire [63:0] zext_ln529_fu_1225_p1;
  reg [63:0] zext_ln529_reg_1472;
  wire [63:0] zext_ln530_fu_1236_p1;
  reg [63:0] zext_ln530_reg_1482;
  wire [63:0] zext_ln531_fu_1246_p1;
  reg [63:0] zext_ln531_reg_1492;
  wire ap_CS_fsm_state13;
  wire [63:0] zext_ln532_fu_1256_p1;
  reg [63:0] zext_ln532_reg_1502;
  reg [4:0] ret_address0;
  reg ret_ce0;
  reg ret_we0;
  wire [31:0] ret_q0;
  reg [4:0] ret_address1;
  reg ret_ce1;
  wire [31:0] ret_q1;
  reg [2:0] j_0_reg_276;
  wire ap_CS_fsm_state5;
  reg [2:0] j_assign_reg_287;
  reg [2:0] i_assign_reg_298;
  wire ap_CS_fsm_state11;
  reg [2:0] i_1_reg_309;
  wire ap_CS_fsm_state14;
  wire [63:0] zext_ln511_1_fu_391_p1;
  wire [63:0] zext_ln512_1_fu_406_p1;
  wire [63:0] zext_ln511_fu_423_p1;
  wire [63:0] zext_ln512_fu_434_p1;
  wire [63:0] zext_ln513_1_fu_448_p1;
  wire [63:0] zext_ln514_1_fu_459_p1;
  wire [63:0] zext_ln513_fu_469_p1;
  wire [63:0] zext_ln514_fu_479_p1;
  wire [63:0] zext_ln457_fu_551_p1;
  wire [63:0] zext_ln473_fu_652_p1;
  wire [63:0] zext_ln486_fu_669_p1;
  wire [5:0] zext_ln508_fu_370_p1;
  wire [7:0] zext_ln511_3_fu_396_p1;
  wire [7:0] add_ln512_fu_400_p2;
  wire [1:0] trunc_ln511_fu_411_p1;
  wire [3:0] or_ln512_fu_428_p2;
  wire [8:0] zext_ln511_2_fu_439_p1;
  wire [8:0] add_ln513_fu_442_p2;
  wire [8:0] add_ln514_fu_453_p2;
  wire [3:0] or_ln513_fu_464_p2;
  wire [3:0] or_ln514_fu_474_p2;
  wire [3:0] zext_ln517_fu_508_p1;
  wire [3:0] add_ln444_fu_524_p2;
  wire [1:0] add_ln457_1_fu_538_p2;
  wire [3:0] or_ln_fu_544_p3;
  wire [23:0] grp_fu_332_p4;
  wire [31:0] and_ln_fu_556_p3;
  wire [23:0] grp_fu_342_p4;
  wire [31:0] and_ln3_fu_578_p3;
  wire [29:0] trunc_ln459_fu_592_p1;
  wire [30:0] tmp_fu_596_p3;
  wire [29:0] trunc_ln460_fu_610_p1;
  wire [0:0] icmp_ln458_fu_586_p2;
  wire [30:0] xor_ln460_fu_604_p2;
  wire [30:0] tmp_1_fu_614_p3;
  wire [1:0] xor_ln473_fu_640_p2;
  wire [3:0] or_ln1_fu_645_p3;
  wire [1:0] add_ln486_fu_657_p2;
  wire [3:0] or_ln2_fu_662_p3;
  wire [30:0] trunc_ln_fu_674_p3;
  wire [30:0] xor_ln445_fu_681_p2;
  wire [30:0] select_ln445_fu_687_p3;
  wire [30:0] xor_ln448_fu_694_p2;
  wire [23:0] tmp_6_fu_699_p4;
  wire [31:0] and_ln1_fu_709_p3;
  wire [30:0] shl_ln450_fu_723_p2;
  wire [0:0] icmp_ln449_fu_717_p2;
  wire [30:0] xor_ln449_fu_729_p2;
  wire [30:0] select_ln449_fu_735_p3;
  wire [30:0] xor_ln452_fu_743_p2;
  wire [23:0] tmp_8_fu_756_p4;
  wire [31:0] and_ln2_fu_766_p3;
  wire [31:0] x_assign_2_fu_748_p3;
  wire [0:0] icmp_ln453_fu_774_p2;
  wire [31:0] xor_ln454_fu_780_p2;
  wire [31:0] and_ln4_fu_797_p3;
  wire [30:0] shl_ln462_fu_810_p2;
  wire [0:0] icmp_ln461_fu_804_p2;
  wire [30:0] xor_ln461_fu_815_p2;
  wire [30:0] select_ln461_fu_821_p3;
  wire [30:0] trunc_ln457_1_fu_794_p1;
  wire [30:0] xor_ln464_fu_829_p2;
  wire [23:0] tmp_3_fu_843_p4;
  wire [31:0] and_ln5_fu_853_p3;
  wire [31:0] x_assign_9_fu_835_p3;
  wire [0:0] icmp_ln465_fu_861_p2;
  wire [31:0] xor_ln466_fu_867_p2;
  wire [31:0] and_ln6_fu_881_p3;
  wire [29:0] trunc_ln475_fu_895_p1;
  wire [30:0] trunc_ln6_fu_899_p3;
  wire [0:0] icmp_ln474_fu_889_p2;
  wire [30:0] xor_ln474_fu_907_p2;
  wire [30:0] select_ln474_fu_913_p3;
  wire [30:0] trunc_ln476_fu_921_p1;
  wire [31:0] and_ln9_fu_941_p3;
  wire [29:0] trunc_ln488_fu_955_p1;
  wire [30:0] tmp_11_fu_959_p3;
  wire [29:0] trunc_ln489_fu_973_p1;
  wire [0:0] icmp_ln487_fu_949_p2;
  wire [30:0] xor_ln489_fu_967_p2;
  wire [30:0] tmp_12_fu_977_p3;
  wire [31:0] select_ln465_fu_873_p3;
  wire [31:0] select_ln453_fu_786_p3;
  wire [31:0] and_ln7_fu_1009_p3;
  wire [30:0] shl_ln479_fu_1022_p2;
  wire [0:0] icmp_ln478_fu_1016_p2;
  wire [30:0] xor_ln480_fu_1027_p2;
  wire [30:0] shl_ln480_fu_1033_p2;
  wire [30:0] select_ln478_fu_1038_p3;
  wire [23:0] tmp_9_fu_1054_p4;
  wire [31:0] and_ln8_fu_1064_p3;
  wire [31:0] x_assign_1_fu_1046_p3;
  wire [0:0] icmp_ln481_fu_1072_p2;
  wire [31:0] xor_ln482_fu_1078_p2;
  wire [31:0] and_ln10_fu_1092_p3;
  wire [30:0] shl_ln491_fu_1105_p2;
  wire [0:0] icmp_ln490_fu_1099_p2;
  wire [30:0] xor_ln492_fu_1110_p2;
  wire [30:0] shl_ln492_fu_1116_p2;
  wire [30:0] select_ln490_fu_1121_p3;
  wire [23:0] tmp_14_fu_1137_p4;
  wire [31:0] and_ln11_fu_1147_p3;
  wire [31:0] x_assign_6_fu_1129_p3;
  wire [0:0] icmp_ln493_fu_1155_p2;
  wire [31:0] xor_ln494_fu_1161_p2;
  wire [31:0] xor_ln524_1_fu_1175_p2;
  wire [31:0] select_ln481_fu_1084_p3;
  wire [31:0] select_ln493_fu_1167_p3;
  wire [31:0] xor_ln524_4_fu_1184_p2;
  wire [31:0] xor_ln524_5_fu_1190_p2;
  wire [31:0] xor_ln524_2_fu_1179_p2;
  wire [1:0] trunc_ln529_fu_1213_p1;
  wire [3:0] or_ln530_fu_1230_p2;
  wire [3:0] or_ln531_fu_1241_p2;
  wire [3:0] or_ln532_fu_1251_p2;
  reg [13:0] ap_NS_fsm;

  initial begin
    #0 ap_CS_fsm = 14'd1;
  end


  AddRoundKey_Invercud
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  ret_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ret_address0),
    .ce0(ret_ce0),
    .we0(ret_we0),
    .d0(xor_ln524_reg_1453),
    .q0(ret_q0),
    .address1(ret_address1),
    .ce1(ret_ce1),
    .q1(ret_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state6) & (icmp_ln516_fu_484_p2 == 1'd1)) begin
      i_1_reg_309 <= 3'd0;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      i_1_reg_309 <= i_reg_1461;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln516_fu_484_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      i_assign_reg_298 <= 3'd0;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      i_assign_reg_298 <= i_3_reg_1348;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      j_0_reg_276 <= j_reg_1269;
    end else if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      j_0_reg_276 <= 3'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln508_fu_374_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      j_assign_reg_287 <= 3'd0;
    end else if((1'b1 == ap_CS_fsm_state7) & (icmp_ln517_fu_512_p2 == 1'd1)) begin
      j_assign_reg_287 <= j_1_reg_1328;
    end 
  end

  assign shl_ln_fu_415_p3_temp_3 = shl_ln_fu_415_p3 & 3'd12;
  assign shl_ln_reg_1289_temp_4 = shl_ln_reg_1289 & 3'd3;
  assign shl_ln_fu_415_p3_temp_3_temp_5 = shl_ln_fu_415_p3_temp_3 | shl_ln_reg_1289_temp_4;
  assign zext_ln512_fu_434_p1_temp_6 = zext_ln512_fu_434_p1 & 63'd12;
  assign statemt_addr_16_reg_1300_temp_7 = statemt_addr_16_reg_1300 & 4'd19;
  assign zext_ln512_fu_434_p1_temp_6_temp_8 = zext_ln512_fu_434_p1_temp_6 | statemt_addr_16_reg_1300_temp_7;
  assign zext_ln511_fu_423_p1_temp_9 = zext_ln511_fu_423_p1 & 63'd12;
  assign statemt_addr_reg_1295_temp_10 = statemt_addr_reg_1295 & 4'd19;
  assign zext_ln511_fu_423_p1_temp_9_temp_11 = zext_ln511_fu_423_p1_temp_9 | statemt_addr_reg_1295_temp_10;

  always @(posedge ap_clk) begin
    if((icmp_ln508_fu_374_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      add_ln511_reg_1274 <= add_ln511_fu_386_p2;
      shl_ln_reg_1289 <= shl_ln_fu_415_p3_temp_3_temp_5;
      statemt_addr_16_reg_1300 <= zext_ln512_fu_434_p1_temp_6_temp_8;
      statemt_addr_reg_1295 <= zext_ln511_fu_423_p1_temp_9_temp_11;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      i_3_reg_1348 <= i_3_fu_518_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      i_reg_1461 <= i_fu_1207_p2;
    end 
  end

  assign select_ln458_fu_622_p3_temp_12 = select_ln458_fu_622_p3 >> 1'd7;
  assign select_ln458_fu_622_p3_temp_13 = select_ln458_fu_622_p3_temp_12 & 24'd16777215;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      icmp_ln445_reg_1374 <= icmp_ln445_fu_564_p2;
      select_ln458_reg_1396 <= select_ln458_fu_622_p3;
      statemt_load_33_reg_1390 <= statemt_q1;
      tmp_2_reg_1401 <= select_ln458_fu_622_p3_temp_13;
      trunc_ln446_reg_1379 <= trunc_ln446_fu_570_p1;
      trunc_ln447_reg_1384 <= trunc_ln447_fu_574_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      j_1_reg_1328 <= j_1_fu_490_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      j_reg_1269 <= j_fu_380_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3)) begin
      reg_352 <= grp_fu_320_p2;
      reg_357 <= grp_fu_326_p2;
    end 
  end

  assign select_ln487_fu_985_p3_temp_14 = select_ln487_fu_985_p3 >> 1'd7;
  assign select_ln487_fu_985_p3_temp_15 = select_ln487_fu_985_p3_temp_14 & 24'd16777215;
  assign xor_ln477_fu_925_p2_temp_16 = xor_ln477_fu_925_p2 >> 1'd7;
  assign xor_ln477_fu_925_p2_temp_17 = xor_ln477_fu_925_p2_temp_16 & 24'd16777215;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      select_ln487_reg_1437 <= select_ln487_fu_985_p3;
      statemt_load_34_reg_1416 <= statemt_q0;
      statemt_load_35_reg_1432 <= statemt_q1;
      tmp_13_reg_1443 <= select_ln487_fu_985_p3_temp_15;
      tmp_7_reg_1427 <= xor_ln477_fu_925_p2_temp_17;
      xor_ln477_reg_1421 <= xor_ln477_fu_925_p2;
      xor_ln524_3_reg_1448 <= xor_ln524_3_fu_1003_p2;
    end 
  end

  assign shl_ln1_fu_500_p3_temp_18 = shl_ln1_fu_500_p3 & 3'd12;
  assign shl_ln1_reg_1340_temp_19 = shl_ln1_reg_1340 & 3'd3;
  assign shl_ln1_fu_500_p3_temp_18_temp_20 = shl_ln1_fu_500_p3_temp_18 | shl_ln1_reg_1340_temp_19;

  always @(posedge ap_clk) begin
    if((icmp_ln516_fu_484_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      shl_ln1_reg_1340 <= shl_ln1_fu_500_p3_temp_18_temp_20;
      trunc_ln521_reg_1333 <= trunc_ln521_fu_496_p1;
    end 
  end

  assign shl_ln2_fu_1217_p3_temp_21 = shl_ln2_fu_1217_p3 & 3'd12;
  assign shl_ln2_reg_1466_temp_22 = shl_ln2_reg_1466 & 3'd3;
  assign shl_ln2_fu_1217_p3_temp_21_temp_23 = shl_ln2_fu_1217_p3_temp_21 | shl_ln2_reg_1466_temp_22;
  assign zext_ln529_fu_1225_p1_temp_24 = zext_ln529_fu_1225_p1 & 63'd12;
  assign zext_ln529_reg_1472_temp_25 = zext_ln529_reg_1472 & 63'd18446744073709551603;
  assign zext_ln529_fu_1225_p1_temp_24_temp_26 = zext_ln529_fu_1225_p1_temp_24 | zext_ln529_reg_1472_temp_25;
  assign zext_ln530_fu_1236_p1_temp_27 = zext_ln530_fu_1236_p1 & 63'd12;
  assign zext_ln530_reg_1482_temp_28 = zext_ln530_reg_1482 & 63'd18446744073709551603;
  assign zext_ln530_fu_1236_p1_temp_27_temp_29 = zext_ln530_fu_1236_p1_temp_27 | zext_ln530_reg_1482_temp_28;

  always @(posedge ap_clk) begin
    if((icmp_ln527_fu_1201_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state12)) begin
      shl_ln2_reg_1466 <= shl_ln2_fu_1217_p3_temp_21_temp_23;
      zext_ln529_reg_1472 <= zext_ln529_fu_1225_p1_temp_24_temp_26;
      zext_ln530_reg_1482 <= zext_ln530_fu_1236_p1_temp_27_temp_29;
    end 
  end

  assign shl_ln511_1_fu_362_p3_temp_30 = shl_ln511_1_fu_362_p3 & 5'd60;
  assign shl_ln511_1_reg_1261_temp_31 = shl_ln511_1_reg_1261 & 5'd3;
  assign shl_ln511_1_fu_362_p3_temp_30_temp_32 = shl_ln511_1_fu_362_p3_temp_30 | shl_ln511_1_reg_1261_temp_31;

  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
      shl_ln511_1_reg_1261 <= shl_ln511_1_fu_362_p3_temp_30_temp_32;
    end 
  end

  assign zext_ln513_fu_469_p1_temp_33 = zext_ln513_fu_469_p1 & 63'd12;
  assign statemt_addr_17_reg_1315_temp_34 = statemt_addr_17_reg_1315 & 4'd19;
  assign zext_ln513_fu_469_p1_temp_33_temp_35 = zext_ln513_fu_469_p1_temp_33 | statemt_addr_17_reg_1315_temp_34;
  assign zext_ln514_fu_479_p1_temp_36 = zext_ln514_fu_479_p1 & 63'd12;
  assign statemt_addr_18_reg_1320_temp_37 = statemt_addr_18_reg_1320 & 4'd19;
  assign zext_ln514_fu_479_p1_temp_36_temp_38 = zext_ln514_fu_479_p1_temp_36 | statemt_addr_18_reg_1320_temp_37;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_addr_17_reg_1315 <= zext_ln513_fu_469_p1_temp_33_temp_35;
      statemt_addr_18_reg_1320 <= zext_ln514_fu_479_p1_temp_36_temp_38;
    end 
  end

  assign zext_ln444_fu_529_p1_temp_39 = zext_ln444_fu_529_p1 & 4'd15;
  assign zext_ln444_reg_1353_temp_40 = zext_ln444_reg_1353 & 4'd18446744073709551600;
  assign zext_ln444_fu_529_p1_temp_39_temp_41 = zext_ln444_fu_529_p1_temp_39 | zext_ln444_reg_1353_temp_40;

  always @(posedge ap_clk) begin
    if((icmp_ln517_fu_512_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      trunc_ln457_reg_1363 <= trunc_ln457_fu_534_p1;
      zext_ln444_reg_1353 <= zext_ln444_fu_529_p1_temp_39_temp_41;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      xor_ln524_reg_1453 <= xor_ln524_fu_1195_p2;
    end 
  end

  assign zext_ln531_fu_1246_p1_temp_42 = zext_ln531_fu_1246_p1 & 63'd12;
  assign zext_ln531_reg_1492_temp_43 = zext_ln531_reg_1492 & 63'd18446744073709551603;
  assign zext_ln531_fu_1246_p1_temp_42_temp_44 = zext_ln531_fu_1246_p1_temp_42 | zext_ln531_reg_1492_temp_43;
  assign zext_ln532_fu_1256_p1_temp_45 = zext_ln532_fu_1256_p1 & 63'd12;
  assign zext_ln532_reg_1502_temp_46 = zext_ln532_reg_1502 & 63'd18446744073709551603;
  assign zext_ln532_fu_1256_p1_temp_45_temp_47 = zext_ln532_fu_1256_p1_temp_45 | zext_ln532_reg_1502_temp_46;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      zext_ln531_reg_1492 <= zext_ln531_fu_1246_p1_temp_42_temp_44;
      zext_ln532_reg_1502 <= zext_ln532_fu_1256_p1_temp_45_temp_47;
    end 
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1) | (1'b1 == ap_CS_fsm_state12) & (icmp_ln527_fu_1201_p2 == 1'd1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state12) & (icmp_ln527_fu_1201_p2 == 1'd1)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      ret_address0 = zext_ln532_fu_1256_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      ret_address0 = zext_ln529_fu_1225_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      ret_address0 = zext_ln444_reg_1353;
    end else begin
      ret_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      ret_address1 = zext_ln531_fu_1246_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      ret_address1 = zext_ln530_fu_1236_p1;
    end else begin
      ret_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12)) begin
      ret_ce0 = 1'b1;
    end else begin
      ret_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12)) begin
      ret_ce1 = 1'b1;
    end else begin
      ret_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      ret_we0 = 1'b1;
    end else begin
      ret_we0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address0 = zext_ln531_reg_1492;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address0 = zext_ln529_reg_1472;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = zext_ln473_fu_652_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address0 = zext_ln444_fu_529_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address0 = statemt_addr_17_reg_1315;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address0 = statemt_addr_reg_1295;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = zext_ln513_fu_469_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address0 = zext_ln511_fu_423_p1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address1 = zext_ln532_reg_1502;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address1 = zext_ln530_reg_1482;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = zext_ln486_fu_669_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address1 = zext_ln457_fu_551_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address1 = statemt_addr_18_reg_1320;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address1 = statemt_addr_16_reg_1300;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address1 = zext_ln514_fu_479_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address1 = zext_ln512_fu_434_p1;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state7)) begin
      statemt_ce1 = 1'b1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d0 = ret_q1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d0 = ret_q0;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d0 = reg_352;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d1 = ret_q0;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d1 = ret_q1;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d1 = reg_357;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt_we1 = 1'b1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address0 = zext_ln513_1_fu_448_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address0 = zext_ln511_1_fu_391_p1;
    end else begin
      word_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address1 = zext_ln514_1_fu_459_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address1 = zext_ln512_1_fu_406_p1;
    end else begin
      word_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce0 = 1'b1;
    end else begin
      word_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce1 = 1'b1;
    end else begin
      word_ce1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((icmp_ln508_fu_374_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state6: begin
        if((1'b1 == ap_CS_fsm_state6) & (icmp_ln516_fu_484_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end
      end
      ap_ST_fsm_state7: begin
        if((1'b1 == ap_CS_fsm_state7) & (icmp_ln517_fu_512_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state12: begin
        if((1'b1 == ap_CS_fsm_state12) & (icmp_ln527_fu_1201_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state13;
        end
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign add_ln444_fu_524_p2 = zext_ln517_fu_508_p1 + shl_ln1_reg_1340;
  assign add_ln457_1_fu_538_p2 = trunc_ln457_fu_534_p1 + 2'd1;
  assign add_ln486_fu_657_p2 = $signed(trunc_ln457_reg_1363) + $signed(2'd3);
  assign add_ln511_fu_386_p2 = zext_ln508_fu_370_p1 + shl_ln511_1_reg_1261;
  assign add_ln512_fu_400_p2 = 8'd120 + zext_ln511_3_fu_396_p1;
  assign add_ln513_fu_442_p2 = 9'd240 + zext_ln511_2_fu_439_p1;
  assign add_ln514_fu_453_p2 = $signed(9'd360) + $signed(zext_ln511_2_fu_439_p1);
  assign tmp_13_reg_1443_temp_48 = tmp_13_reg_1443 << 1'd8;
  assign and_ln10_fu_1092_p3 = tmp_13_reg_1443_temp_48;
  assign tmp_14_fu_1137_p4_temp_49 = tmp_14_fu_1137_p4 << 1'd8;
  assign and_ln11_fu_1147_p3 = tmp_14_fu_1137_p4_temp_49;
  assign tmp_6_fu_699_p4_temp_50 = tmp_6_fu_699_p4 << 1'd8;
  assign and_ln1_fu_709_p3 = tmp_6_fu_699_p4_temp_50;
  assign tmp_8_fu_756_p4_temp_51 = tmp_8_fu_756_p4 << 1'd8;
  assign and_ln2_fu_766_p3 = tmp_8_fu_756_p4_temp_51;
  assign grp_fu_342_p4_temp_52 = grp_fu_342_p4 << 1'd8;
  assign and_ln3_fu_578_p3 = grp_fu_342_p4_temp_52;
  assign tmp_2_reg_1401_temp_53 = tmp_2_reg_1401 << 1'd8;
  assign and_ln4_fu_797_p3 = tmp_2_reg_1401_temp_53;
  assign tmp_3_fu_843_p4_temp_54 = tmp_3_fu_843_p4 << 1'd8;
  assign and_ln5_fu_853_p3 = tmp_3_fu_843_p4_temp_54;
  assign grp_fu_332_p4_temp_55 = grp_fu_332_p4 << 1'd8;
  assign and_ln6_fu_881_p3 = grp_fu_332_p4_temp_55;
  assign tmp_7_reg_1427_temp_56 = tmp_7_reg_1427 << 1'd8;
  assign and_ln7_fu_1009_p3 = tmp_7_reg_1427_temp_56;
  assign tmp_9_fu_1054_p4_temp_57 = tmp_9_fu_1054_p4 << 1'd8;
  assign and_ln8_fu_1064_p3 = tmp_9_fu_1054_p4_temp_57;
  assign grp_fu_342_p4_temp_58 = grp_fu_342_p4 << 1'd8;
  assign and_ln9_fu_941_p3 = grp_fu_342_p4_temp_58;
  assign grp_fu_332_p4_temp_59 = grp_fu_332_p4 << 1'd8;
  assign and_ln_fu_556_p3 = grp_fu_332_p4_temp_59;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign grp_fu_320_p2 = word_q0 ^ statemt_q0;
  assign grp_fu_326_p2 = word_q1 ^ statemt_q1;
  assign statemt_q0_temp_60 = statemt_q0 >> 1'd7;
  assign statemt_q0_temp_61 = statemt_q0_temp_60 & 24'd16777215;
  assign grp_fu_332_p4 = statemt_q0_temp_61;
  assign statemt_q1_temp_62 = statemt_q1 >> 1'd7;
  assign statemt_q1_temp_63 = statemt_q1_temp_62 & 24'd16777215;
  assign grp_fu_342_p4 = statemt_q1_temp_63;
  assign i_3_fu_518_p2 = i_assign_reg_298 + 3'd1;
  assign i_fu_1207_p2 = i_1_reg_309 + 3'd1;
  assign icmp_ln445_fu_564_p2 = (and_ln_fu_556_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln449_fu_717_p2 = (and_ln1_fu_709_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln453_fu_774_p2 = (and_ln2_fu_766_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln458_fu_586_p2 = (and_ln3_fu_578_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln461_fu_804_p2 = (and_ln4_fu_797_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln465_fu_861_p2 = (and_ln5_fu_853_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln474_fu_889_p2 = (and_ln6_fu_881_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln478_fu_1016_p2 = (and_ln7_fu_1009_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln481_fu_1072_p2 = (and_ln8_fu_1064_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln487_fu_949_p2 = (and_ln9_fu_941_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln490_fu_1099_p2 = (and_ln10_fu_1092_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln493_fu_1155_p2 = (and_ln11_fu_1147_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln508_fu_374_p2 = (j_0_reg_276 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln516_fu_484_p2 = (j_assign_reg_287 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln517_fu_512_p2 = (i_assign_reg_298 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln527_fu_1201_p2 = (i_1_reg_309 == 3'd4)? 1'b1 : 1'b0;
  assign j_1_fu_490_p2 = j_assign_reg_287 + 3'd1;
  assign j_fu_380_p2 = j_0_reg_276 + 3'd1;
  assign trunc_ln521_reg_1333_temp_64 = trunc_ln521_reg_1333 << 1'd2;
  assign trunc_ln521_reg_1333_temp_65 = trunc_ln521_reg_1333_temp_64 | xor_ln473_fu_640_p2;
  assign or_ln1_fu_645_p3 = trunc_ln521_reg_1333_temp_65;
  assign trunc_ln521_reg_1333_temp_66 = trunc_ln521_reg_1333 << 1'd2;
  assign trunc_ln521_reg_1333_temp_67 = trunc_ln521_reg_1333_temp_66 | add_ln486_fu_657_p2;
  assign or_ln2_fu_662_p3 = trunc_ln521_reg_1333_temp_67;
  assign or_ln512_fu_428_p2 = shl_ln_fu_415_p3 | 4'd1;
  assign or_ln513_fu_464_p2 = shl_ln_reg_1289 | 4'd2;
  assign or_ln514_fu_474_p2 = shl_ln_reg_1289 | 4'd3;
  assign or_ln530_fu_1230_p2 = shl_ln2_fu_1217_p3 | 4'd1;
  assign or_ln531_fu_1241_p2 = shl_ln2_reg_1466 | 4'd2;
  assign or_ln532_fu_1251_p2 = shl_ln2_reg_1466 | 4'd3;
  assign trunc_ln521_reg_1333_temp_68 = trunc_ln521_reg_1333 << 1'd2;
  assign trunc_ln521_reg_1333_temp_69 = trunc_ln521_reg_1333_temp_68 | add_ln457_1_fu_538_p2;
  assign or_ln_fu_544_p3 = trunc_ln521_reg_1333_temp_69;
  assign icmp_ln445_reg_1374_temp_70 = icmp_ln445_reg_1374 & 30'd1;
  assign select_ln445_fu_687_p3 = (icmp_ln445_reg_1374_temp_70 === 1'b1)? xor_ln445_fu_681_p2 : trunc_ln_fu_674_p3;
  assign icmp_ln449_fu_717_p2_temp_71 = icmp_ln449_fu_717_p2 & 30'd1;
  assign select_ln449_fu_735_p3 = (icmp_ln449_fu_717_p2_temp_71 === 1'b1)? xor_ln449_fu_729_p2 : shl_ln450_fu_723_p2;
  assign icmp_ln453_fu_774_p2_temp_72 = icmp_ln453_fu_774_p2 & 31'd1;
  assign select_ln453_fu_786_p3 = (icmp_ln453_fu_774_p2_temp_72 === 1'b1)? xor_ln454_fu_780_p2 : x_assign_2_fu_748_p3;
  assign icmp_ln458_fu_586_p2_temp_73 = icmp_ln458_fu_586_p2 & 30'd1;
  assign select_ln458_fu_622_p3 = (icmp_ln458_fu_586_p2_temp_73 === 1'b1)? xor_ln460_fu_604_p2 : tmp_1_fu_614_p3;
  assign icmp_ln461_fu_804_p2_temp_74 = icmp_ln461_fu_804_p2 & 30'd1;
  assign select_ln461_fu_821_p3 = (icmp_ln461_fu_804_p2_temp_74 === 1'b1)? xor_ln461_fu_815_p2 : shl_ln462_fu_810_p2;
  assign icmp_ln465_fu_861_p2_temp_75 = icmp_ln465_fu_861_p2 & 31'd1;
  assign select_ln465_fu_873_p3 = (icmp_ln465_fu_861_p2_temp_75 === 1'b1)? xor_ln466_fu_867_p2 : x_assign_9_fu_835_p3;
  assign icmp_ln474_fu_889_p2_temp_76 = icmp_ln474_fu_889_p2 & 30'd1;
  assign select_ln474_fu_913_p3 = (icmp_ln474_fu_889_p2_temp_76 === 1'b1)? xor_ln474_fu_907_p2 : trunc_ln6_fu_899_p3;
  assign icmp_ln478_fu_1016_p2_temp_77 = icmp_ln478_fu_1016_p2 & 30'd1;
  assign select_ln478_fu_1038_p3 = (icmp_ln478_fu_1016_p2_temp_77 === 1'b1)? xor_ln480_fu_1027_p2 : shl_ln480_fu_1033_p2;
  assign icmp_ln481_fu_1072_p2_temp_78 = icmp_ln481_fu_1072_p2 & 31'd1;
  assign select_ln481_fu_1084_p3 = (icmp_ln481_fu_1072_p2_temp_78 === 1'b1)? xor_ln482_fu_1078_p2 : x_assign_1_fu_1046_p3;
  assign icmp_ln487_fu_949_p2_temp_79 = icmp_ln487_fu_949_p2 & 30'd1;
  assign select_ln487_fu_985_p3 = (icmp_ln487_fu_949_p2_temp_79 === 1'b1)? xor_ln489_fu_967_p2 : tmp_12_fu_977_p3;
  assign icmp_ln490_fu_1099_p2_temp_80 = icmp_ln490_fu_1099_p2 & 30'd1;
  assign select_ln490_fu_1121_p3 = (icmp_ln490_fu_1099_p2_temp_80 === 1'b1)? xor_ln492_fu_1110_p2 : shl_ln492_fu_1116_p2;
  assign icmp_ln493_fu_1155_p2_temp_81 = icmp_ln493_fu_1155_p2 & 31'd1;
  assign select_ln493_fu_1167_p3 = (icmp_ln493_fu_1155_p2_temp_81 === 1'b1)? xor_ln494_fu_1161_p2 : x_assign_6_fu_1129_p3;
  assign trunc_ln521_fu_496_p1_temp_82 = trunc_ln521_fu_496_p1 << 1'd2;
  assign shl_ln1_fu_500_p3 = trunc_ln521_fu_496_p1_temp_82;
  assign trunc_ln529_fu_1213_p1_temp_83 = trunc_ln529_fu_1213_p1 << 1'd2;
  assign shl_ln2_fu_1217_p3 = trunc_ln529_fu_1213_p1_temp_83;
  assign shl_ln450_fu_723_p2 = xor_ln448_fu_694_p2 << 31'd1;
  assign shl_ln462_fu_810_p2 = select_ln458_reg_1396 << 31'd1;
  assign shl_ln479_fu_1022_p2 = xor_ln477_reg_1421 << 31'd1;
  assign shl_ln480_fu_1033_p2 = xor_ln477_reg_1421 << 31'd1;
  assign shl_ln491_fu_1105_p2 = select_ln487_reg_1437 << 31'd1;
  assign shl_ln492_fu_1116_p2 = select_ln487_reg_1437 << 31'd1;
  assign n_temp_84 = n << 1'd2;
  assign shl_ln511_1_fu_362_p3 = n_temp_84;
  assign trunc_ln511_fu_411_p1_temp_85 = trunc_ln511_fu_411_p1 << 1'd2;
  assign shl_ln_fu_415_p3 = trunc_ln511_fu_411_p1_temp_85;
  assign trunc_ln488_fu_955_p1_temp_86 = trunc_ln488_fu_955_p1 << 1'd1;
  assign tmp_11_fu_959_p3 = trunc_ln488_fu_955_p1_temp_86;
  assign trunc_ln489_fu_973_p1_temp_87 = trunc_ln489_fu_973_p1 << 1'd1;
  assign tmp_12_fu_977_p3 = trunc_ln489_fu_973_p1_temp_87;
  assign select_ln490_fu_1121_p3_temp_88 = select_ln490_fu_1121_p3 >> 1'd7;
  assign select_ln490_fu_1121_p3_temp_89 = select_ln490_fu_1121_p3_temp_88 & 24'd16777215;
  assign tmp_14_fu_1137_p4 = select_ln490_fu_1121_p3_temp_89;
  assign trunc_ln460_fu_610_p1_temp_90 = trunc_ln460_fu_610_p1 << 1'd1;
  assign tmp_1_fu_614_p3 = trunc_ln460_fu_610_p1_temp_90;
  assign xor_ln464_fu_829_p2_temp_91 = xor_ln464_fu_829_p2 >> 1'd7;
  assign xor_ln464_fu_829_p2_temp_92 = xor_ln464_fu_829_p2_temp_91 & 24'd16777215;
  assign tmp_3_fu_843_p4 = xor_ln464_fu_829_p2_temp_92;
  assign xor_ln448_fu_694_p2_temp_93 = xor_ln448_fu_694_p2 >> 1'd7;
  assign xor_ln448_fu_694_p2_temp_94 = xor_ln448_fu_694_p2_temp_93 & 24'd16777215;
  assign tmp_6_fu_699_p4 = xor_ln448_fu_694_p2_temp_94;
  assign xor_ln452_fu_743_p2_temp_95 = xor_ln452_fu_743_p2 >> 1'd7;
  assign xor_ln452_fu_743_p2_temp_96 = xor_ln452_fu_743_p2_temp_95 & 24'd16777215;
  assign tmp_8_fu_756_p4 = xor_ln452_fu_743_p2_temp_96;
  assign select_ln478_fu_1038_p3_temp_97 = select_ln478_fu_1038_p3 >> 1'd7;
  assign select_ln478_fu_1038_p3_temp_98 = select_ln478_fu_1038_p3_temp_97 & 24'd16777215;
  assign tmp_9_fu_1054_p4 = select_ln478_fu_1038_p3_temp_98;
  assign trunc_ln459_fu_592_p1_temp_99 = trunc_ln459_fu_592_p1 << 1'd1;
  assign tmp_fu_596_p3 = trunc_ln459_fu_592_p1_temp_99;
  assign trunc_ln446_fu_570_p1 = (statemt_q0 & 30'd1073741823);
  assign trunc_ln447_fu_574_p1 = (statemt_q0 & 31'd2147483647);
  assign trunc_ln457_1_fu_794_p1 = (statemt_load_33_reg_1390 & 31'd2147483647);
  assign trunc_ln457_fu_534_p1 = (i_assign_reg_298 & 2'd3);
  assign trunc_ln459_fu_592_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln460_fu_610_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln475_fu_895_p1 = (statemt_q0 & 30'd1073741823);
  assign trunc_ln476_fu_921_p1 = (statemt_q0 & 31'd2147483647);
  assign trunc_ln488_fu_955_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln489_fu_973_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln511_fu_411_p1 = (j_0_reg_276 & 2'd3);
  assign trunc_ln521_fu_496_p1 = (j_assign_reg_287 & 2'd3);
  assign trunc_ln529_fu_1213_p1 = (i_1_reg_309 & 2'd3);
  assign trunc_ln475_fu_895_p1_temp_100 = trunc_ln475_fu_895_p1 << 1'd1;
  assign trunc_ln6_fu_899_p3 = trunc_ln475_fu_895_p1_temp_100;
  assign trunc_ln446_reg_1379_temp_101 = trunc_ln446_reg_1379 << 1'd1;
  assign trunc_ln_fu_674_p3 = trunc_ln446_reg_1379_temp_101;
  assign select_ln478_fu_1038_p3_temp_102 = select_ln478_fu_1038_p3 << 1'd1;
  assign x_assign_1_fu_1046_p3 = select_ln478_fu_1038_p3_temp_102;
  assign xor_ln452_fu_743_p2_temp_103 = xor_ln452_fu_743_p2 << 1'd1;
  assign x_assign_2_fu_748_p3 = xor_ln452_fu_743_p2_temp_103;
  assign select_ln490_fu_1121_p3_temp_104 = select_ln490_fu_1121_p3 << 1'd1;
  assign x_assign_6_fu_1129_p3 = select_ln490_fu_1121_p3_temp_104;
  assign xor_ln464_fu_829_p2_temp_105 = xor_ln464_fu_829_p2 << 1'd1;
  assign x_assign_9_fu_835_p3 = xor_ln464_fu_829_p2_temp_105;
  assign xor_ln445_fu_681_p2 = trunc_ln_fu_674_p3 ^ 31'd283;
  assign xor_ln448_fu_694_p2 = trunc_ln447_reg_1384 ^ select_ln445_fu_687_p3;
  assign xor_ln449_fu_729_p2 = shl_ln450_fu_723_p2 ^ 31'd283;
  assign xor_ln452_fu_743_p2 = trunc_ln447_reg_1384 ^ select_ln449_fu_735_p3;
  assign xor_ln454_fu_780_p2 = x_assign_2_fu_748_p3 ^ 32'd283;
  assign xor_ln460_fu_604_p2 = tmp_fu_596_p3 ^ 31'd283;
  assign xor_ln461_fu_815_p2 = shl_ln462_fu_810_p2 ^ 31'd283;
  assign xor_ln464_fu_829_p2 = trunc_ln457_1_fu_794_p1 ^ select_ln461_fu_821_p3;
  assign xor_ln466_fu_867_p2 = x_assign_9_fu_835_p3 ^ 32'd283;
  assign xor_ln473_fu_640_p2 = trunc_ln457_reg_1363 ^ 2'd2;
  assign xor_ln474_fu_907_p2 = trunc_ln6_fu_899_p3 ^ 31'd283;
  assign xor_ln477_fu_925_p2 = trunc_ln476_fu_921_p1 ^ select_ln474_fu_913_p3;
  assign xor_ln480_fu_1027_p2 = shl_ln479_fu_1022_p2 ^ 31'd283;
  assign xor_ln482_fu_1078_p2 = x_assign_1_fu_1046_p3 ^ 32'd283;
  assign xor_ln489_fu_967_p2 = tmp_11_fu_959_p3 ^ 31'd283;
  assign xor_ln492_fu_1110_p2 = shl_ln491_fu_1105_p2 ^ 31'd283;
  assign xor_ln494_fu_1161_p2 = x_assign_6_fu_1129_p3 ^ 32'd283;
  assign xor_ln524_1_fu_1175_p2 = statemt_load_35_reg_1432 ^ statemt_load_34_reg_1416;
  assign xor_ln524_2_fu_1179_p2 = xor_ln524_1_fu_1175_p2 ^ statemt_load_33_reg_1390;
  assign xor_ln524_3_fu_1003_p2 = select_ln465_fu_873_p3 ^ select_ln453_fu_786_p3;
  assign xor_ln524_4_fu_1184_p2 = select_ln493_fu_1167_p3 ^ select_ln481_fu_1084_p3;
  assign xor_ln524_5_fu_1190_p2 = xor_ln524_4_fu_1184_p2 ^ xor_ln524_3_reg_1448;
  assign xor_ln524_fu_1195_p2 = xor_ln524_5_fu_1190_p2 ^ xor_ln524_2_fu_1179_p2;
  assign zext_ln444_fu_529_p1 = add_ln444_fu_524_p2;
  assign zext_ln457_fu_551_p1 = or_ln_fu_544_p3;
  assign zext_ln473_fu_652_p1 = or_ln1_fu_645_p3;
  assign zext_ln486_fu_669_p1 = or_ln2_fu_662_p3;
  assign zext_ln508_fu_370_p1 = j_0_reg_276;
  assign zext_ln511_1_fu_391_p1 = add_ln511_fu_386_p2;
  assign zext_ln511_2_fu_439_p1 = add_ln511_reg_1274;
  assign zext_ln511_3_fu_396_p1 = add_ln511_fu_386_p2;
  assign zext_ln511_fu_423_p1 = shl_ln_fu_415_p3;
  assign zext_ln512_1_fu_406_p1 = add_ln512_fu_400_p2;
  assign zext_ln512_fu_434_p1 = or_ln512_fu_428_p2;
  assign zext_ln513_1_fu_448_p1 = add_ln513_fu_442_p2;
  assign zext_ln513_fu_469_p1 = or_ln513_fu_464_p2;
  assign zext_ln514_1_fu_459_p1 = add_ln514_fu_453_p2;
  assign zext_ln514_fu_479_p1 = or_ln514_fu_474_p2;
  assign zext_ln517_fu_508_p1 = i_assign_reg_298;
  assign zext_ln529_fu_1225_p1 = shl_ln2_fu_1217_p3;
  assign zext_ln530_fu_1236_p1 = or_ln530_fu_1230_p2;
  assign zext_ln531_fu_1246_p1 = or_ln531_fu_1241_p2;
  assign zext_ln532_fu_1256_p1 = or_ln532_fu_1251_p2;

  always @(posedge ap_clk) begin
    shl_ln511_1_reg_1261 <= shl_ln511_1_reg_1261 & 1'd60;
    shl_ln_reg_1289 <= shl_ln_reg_1289 & 1'd12;
    statemt_addr_reg_1295 <= statemt_addr_reg_1295 & 1'd28;
    statemt_addr_reg_1295 <= statemt_addr_reg_1295 & 4'd15;
    statemt_addr_16_reg_1300 <= statemt_addr_16_reg_1300 & 1'd29;
    statemt_addr_16_reg_1300 <= statemt_addr_16_reg_1300 & 4'd15;
    statemt_addr_17_reg_1315 <= statemt_addr_17_reg_1315 & 1'd30;
    statemt_addr_17_reg_1315 <= statemt_addr_17_reg_1315 & 4'd15;
    statemt_addr_18_reg_1320 <= statemt_addr_18_reg_1320 & 1'd31;
    statemt_addr_18_reg_1320 <= statemt_addr_18_reg_1320 & 4'd15;
    shl_ln1_reg_1340 <= shl_ln1_reg_1340 & 1'd12;
    zext_ln444_reg_1353 <= zext_ln444_reg_1353 & 63'd15;
    shl_ln2_reg_1466 <= shl_ln2_reg_1466 & 1'd12;
    zext_ln529_reg_1472 <= zext_ln529_reg_1472 & 1'd18446744073709551612;
    zext_ln529_reg_1472 <= zext_ln529_reg_1472 & 63'd15;
    zext_ln530_reg_1482 <= zext_ln530_reg_1482 & 1'd18446744073709551613;
    zext_ln530_reg_1482 <= zext_ln530_reg_1482 & 63'd15;
    zext_ln531_reg_1492 <= zext_ln531_reg_1492 & 1'd18446744073709551614;
    zext_ln531_reg_1492 <= zext_ln531_reg_1492 & 63'd15;
    zext_ln532_reg_1502 <= zext_ln532_reg_1502 & 1'd18446744073709551615;
    zext_ln532_reg_1502 <= zext_ln532_reg_1502 & 63'd15;
  end


endmodule

