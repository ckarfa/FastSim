
module AddRoundKey_InversMi
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  statemt_address1,
  statemt_ce1,
  statemt_we1,
  statemt_d1,
  statemt_q1,
  n,
  word_address0,
  word_ce0,
  word_q0,
  word_address1,
  word_ce1,
  word_q1
);

  parameter ap_ST_fsm_state1 = 15'd1;
  parameter ap_ST_fsm_state2 = 15'd2;
  parameter ap_ST_fsm_state3 = 15'd4;
  parameter ap_ST_fsm_state4 = 15'd8;
  parameter ap_ST_fsm_state5 = 15'd16;
  parameter ap_ST_fsm_state6 = 15'd32;
  parameter ap_ST_fsm_state7 = 15'd64;
  parameter ap_ST_fsm_state8 = 15'd128;
  parameter ap_ST_fsm_state9 = 15'd256;
  parameter ap_ST_fsm_state10 = 15'd512;
  parameter ap_ST_fsm_state11 = 15'd1024;
  parameter ap_ST_fsm_state12 = 15'd2048;
  parameter ap_ST_fsm_pp1_stage0 = 15'd4096;
  parameter ap_ST_fsm_pp1_stage1 = 15'd8192;
  parameter ap_ST_fsm_state16 = 15'd16384;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] statemt_address1;
  output statemt_ce1;
  output statemt_we1;
  output [31:0] statemt_d1;
  input [31:0] statemt_q1;
  input [3:0] n;
  output [8:0] word_address0;
  output word_ce0;
  input [31:0] word_q0;
  output [8:0] word_address1;
  output word_ce1;
  input [31:0] word_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  reg [8:0] word_address0;
  reg word_ce0;
  reg [8:0] word_address1;
  reg word_ce1;
  reg [14:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [2:0] i_1_reg_325;
  wire [31:0] grp_fu_336_p2;
  reg [31:0] reg_368;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state4;
  wire [31:0] grp_fu_342_p2;
  reg [31:0] reg_373;
  wire [5:0] shl_ln510_1_fu_378_p3;
  reg [5:0] shl_ln510_1_reg_1277;
  wire [2:0] j_fu_392_p2;
  reg [2:0] j_reg_1285;
  wire ap_CS_fsm_state2;
  wire [5:0] add_ln510_fu_402_p2;
  reg [5:0] add_ln510_reg_1290;
  wire [0:0] icmp_ln507_fu_386_p2;
  wire [3:0] shl_ln_fu_431_p3;
  reg [3:0] shl_ln_reg_1305;
  reg [4:0] statemt_addr_reg_1311;
  reg [4:0] statemt_addr_17_reg_1316;
  reg [4:0] statemt_addr_18_reg_1331;
  reg [4:0] statemt_addr_19_reg_1336;
  wire [0:0] icmp_ln515_fu_500_p2;
  wire ap_CS_fsm_state7;
  wire [2:0] j_1_fu_506_p2;
  reg [2:0] j_1_reg_1345;
  wire [1:0] trunc_ln520_fu_512_p1;
  reg [1:0] trunc_ln520_reg_1350;
  wire [3:0] shl_ln1_fu_516_p3;
  reg [3:0] shl_ln1_reg_1357;
  wire [2:0] i_5_fu_534_p2;
  reg [2:0] i_5_reg_1365;
  wire ap_CS_fsm_state8;
  wire [63:0] zext_ln443_fu_545_p1;
  reg [63:0] zext_ln443_reg_1370;
  wire [0:0] icmp_ln516_fu_528_p2;
  wire [1:0] trunc_ln456_fu_550_p1;
  reg [1:0] trunc_ln456_reg_1380;
  wire [0:0] icmp_ln444_fu_580_p2;
  reg [0:0] icmp_ln444_reg_1391;
  wire ap_CS_fsm_state9;
  wire [29:0] trunc_ln445_fu_586_p1;
  reg [29:0] trunc_ln445_reg_1396;
  wire [30:0] trunc_ln446_fu_590_p1;
  reg [30:0] trunc_ln446_reg_1401;
  reg [31:0] statemt_load_20_reg_1407;
  wire [30:0] select_ln457_fu_638_p3;
  reg [30:0] select_ln457_reg_1413;
  reg [23:0] tmp_5_reg_1418;
  reg [31:0] statemt_load_21_reg_1433;
  wire ap_CS_fsm_state10;
  wire [30:0] xor_ln476_fu_941_p2;
  reg [30:0] xor_ln476_reg_1438;
  reg [23:0] tmp_10_reg_1444;
  reg [31:0] statemt_load_22_reg_1449;
  wire [30:0] select_ln486_fu_1001_p3;
  reg [30:0] select_ln486_reg_1454;
  reg [23:0] tmp_15_reg_1460;
  wire [31:0] xor_ln523_3_fu_1019_p2;
  reg [31:0] xor_ln523_3_reg_1465;
  wire [31:0] xor_ln523_fu_1211_p2;
  reg [31:0] xor_ln523_reg_1470;
  wire ap_CS_fsm_state11;
  wire [0:0] icmp_ln526_fu_1217_p2;
  reg [0:0] icmp_ln526_reg_1475;
  wire ap_CS_fsm_pp1_stage0;
  wire ap_block_state13_pp1_stage0_iter0;
  wire ap_block_state15_pp1_stage0_iter1;
  wire ap_block_pp1_stage0_11001;
  wire [2:0] i_fu_1223_p2;
  reg [2:0] i_reg_1479;
  reg ap_enable_reg_pp1_iter0;
  wire [3:0] shl_ln2_fu_1233_p3;
  reg [3:0] shl_ln2_reg_1484;
  wire [63:0] zext_ln529_fu_1241_p1;
  reg [63:0] zext_ln529_reg_1490;
  wire [63:0] zext_ln530_fu_1252_p1;
  reg [63:0] zext_ln530_reg_1500;
  wire [63:0] zext_ln531_fu_1262_p1;
  reg [63:0] zext_ln531_reg_1510;
  wire ap_CS_fsm_pp1_stage1;
  wire ap_block_state14_pp1_stage1_iter0;
  wire ap_block_pp1_stage1_11001;
  wire [63:0] zext_ln532_fu_1272_p1;
  reg [63:0] zext_ln532_reg_1520;
  wire ap_block_pp1_stage0_subdone;
  reg ap_condition_pp1_exit_iter0_state13;
  reg ap_enable_reg_pp1_iter1;
  wire ap_block_pp1_stage1_subdone;
  reg [4:0] ret_address0;
  reg ret_ce0;
  reg ret_we0;
  wire [31:0] ret_q0;
  reg [4:0] ret_address1;
  reg ret_ce1;
  wire [31:0] ret_q1;
  reg [2:0] j_0_reg_292;
  wire ap_CS_fsm_state5;
  reg [2:0] j_assign_reg_303;
  wire ap_CS_fsm_state6;
  reg [2:0] i_assign_reg_314;
  wire ap_CS_fsm_state12;
  reg [2:0] ap_phi_mux_i_1_phi_fu_329_p4;
  wire ap_block_pp1_stage0;
  wire [63:0] zext_ln510_1_fu_407_p1;
  wire [63:0] zext_ln511_1_fu_422_p1;
  wire [63:0] zext_ln510_fu_439_p1;
  wire [63:0] zext_ln511_fu_450_p1;
  wire [63:0] zext_ln512_1_fu_464_p1;
  wire [63:0] zext_ln513_1_fu_475_p1;
  wire [63:0] zext_ln512_fu_485_p1;
  wire [63:0] zext_ln513_fu_495_p1;
  wire [63:0] zext_ln456_fu_567_p1;
  wire [63:0] zext_ln472_fu_668_p1;
  wire [63:0] zext_ln485_fu_685_p1;
  wire ap_block_pp1_stage1;
  wire [5:0] zext_ln507_fu_398_p1;
  wire [7:0] zext_ln510_3_fu_412_p1;
  wire [7:0] add_ln511_fu_416_p2;
  wire [1:0] trunc_ln510_fu_427_p1;
  wire [3:0] or_ln511_fu_444_p2;
  wire [8:0] zext_ln510_2_fu_455_p1;
  wire [8:0] add_ln512_fu_458_p2;
  wire [8:0] add_ln513_fu_469_p2;
  wire [3:0] or_ln512_fu_480_p2;
  wire [3:0] or_ln513_fu_490_p2;
  wire [3:0] zext_ln516_fu_524_p1;
  wire [3:0] add_ln443_fu_540_p2;
  wire [1:0] add_ln456_1_fu_554_p2;
  wire [3:0] or_ln_fu_560_p3;
  wire [23:0] grp_fu_348_p4;
  wire [31:0] and_ln_fu_572_p3;
  wire [23:0] grp_fu_358_p4;
  wire [31:0] and_ln3_fu_594_p3;
  wire [29:0] trunc_ln458_fu_608_p1;
  wire [30:0] tmp_3_fu_612_p3;
  wire [29:0] trunc_ln459_fu_626_p1;
  wire [0:0] icmp_ln457_fu_602_p2;
  wire [30:0] xor_ln459_fu_620_p2;
  wire [30:0] tmp_4_fu_630_p3;
  wire [1:0] xor_ln472_fu_656_p2;
  wire [3:0] or_ln1_fu_661_p3;
  wire [1:0] add_ln485_fu_673_p2;
  wire [3:0] or_ln2_fu_678_p3;
  wire [30:0] trunc_ln_fu_690_p3;
  wire [30:0] xor_ln444_fu_697_p2;
  wire [30:0] select_ln444_fu_703_p3;
  wire [30:0] xor_ln447_fu_710_p2;
  wire [23:0] tmp_8_fu_715_p4;
  wire [31:0] and_ln1_fu_725_p3;
  wire [30:0] shl_ln449_fu_739_p2;
  wire [0:0] icmp_ln448_fu_733_p2;
  wire [30:0] xor_ln448_fu_745_p2;
  wire [30:0] select_ln448_fu_751_p3;
  wire [30:0] xor_ln451_fu_759_p2;
  wire [23:0] tmp_s_fu_772_p4;
  wire [31:0] and_ln2_fu_782_p3;
  wire [31:0] x_assign_2_fu_764_p3;
  wire [0:0] icmp_ln452_fu_790_p2;
  wire [31:0] xor_ln453_fu_796_p2;
  wire [31:0] and_ln4_fu_813_p3;
  wire [30:0] shl_ln461_fu_826_p2;
  wire [0:0] icmp_ln460_fu_820_p2;
  wire [30:0] xor_ln460_fu_831_p2;
  wire [30:0] select_ln460_fu_837_p3;
  wire [30:0] trunc_ln456_1_fu_810_p1;
  wire [30:0] xor_ln463_fu_845_p2;
  wire [23:0] tmp_7_fu_859_p4;
  wire [31:0] and_ln5_fu_869_p3;
  wire [31:0] x_assign_9_fu_851_p3;
  wire [0:0] icmp_ln464_fu_877_p2;
  wire [31:0] xor_ln465_fu_883_p2;
  wire [31:0] and_ln6_fu_897_p3;
  wire [29:0] trunc_ln474_fu_911_p1;
  wire [30:0] trunc_ln6_fu_915_p3;
  wire [0:0] icmp_ln473_fu_905_p2;
  wire [30:0] xor_ln473_fu_923_p2;
  wire [30:0] select_ln473_fu_929_p3;
  wire [30:0] trunc_ln475_fu_937_p1;
  wire [31:0] and_ln9_fu_957_p3;
  wire [29:0] trunc_ln487_fu_971_p1;
  wire [30:0] tmp_13_fu_975_p3;
  wire [29:0] trunc_ln488_fu_989_p1;
  wire [0:0] icmp_ln486_fu_965_p2;
  wire [30:0] xor_ln488_fu_983_p2;
  wire [30:0] tmp_14_fu_993_p3;
  wire [31:0] select_ln464_fu_889_p3;
  wire [31:0] select_ln452_fu_802_p3;
  wire [31:0] and_ln7_fu_1025_p3;
  wire [30:0] shl_ln478_fu_1038_p2;
  wire [0:0] icmp_ln477_fu_1032_p2;
  wire [30:0] xor_ln479_fu_1043_p2;
  wire [30:0] shl_ln479_fu_1049_p2;
  wire [30:0] select_ln477_fu_1054_p3;
  wire [23:0] tmp_11_fu_1070_p4;
  wire [31:0] and_ln8_fu_1080_p3;
  wire [31:0] x_assign_1_fu_1062_p3;
  wire [0:0] icmp_ln480_fu_1088_p2;
  wire [31:0] xor_ln481_fu_1094_p2;
  wire [31:0] and_ln10_fu_1108_p3;
  wire [30:0] shl_ln490_fu_1121_p2;
  wire [0:0] icmp_ln489_fu_1115_p2;
  wire [30:0] xor_ln491_fu_1126_p2;
  wire [30:0] shl_ln491_fu_1132_p2;
  wire [30:0] select_ln489_fu_1137_p3;
  wire [23:0] tmp_16_fu_1153_p4;
  wire [31:0] and_ln11_fu_1163_p3;
  wire [31:0] x_assign_6_fu_1145_p3;
  wire [0:0] icmp_ln492_fu_1171_p2;
  wire [31:0] xor_ln493_fu_1177_p2;
  wire [31:0] xor_ln523_1_fu_1191_p2;
  wire [31:0] select_ln480_fu_1100_p3;
  wire [31:0] select_ln492_fu_1183_p3;
  wire [31:0] xor_ln523_4_fu_1200_p2;
  wire [31:0] xor_ln523_5_fu_1206_p2;
  wire [31:0] xor_ln523_2_fu_1195_p2;
  wire [1:0] trunc_ln529_fu_1229_p1;
  wire [3:0] or_ln530_fu_1246_p2;
  wire [3:0] or_ln531_fu_1257_p2;
  wire [3:0] or_ln532_fu_1267_p2;
  wire ap_CS_fsm_state16;
  reg [14:0] ap_NS_fsm;
  reg ap_idle_pp1;
  wire ap_enable_pp1;

  initial begin
    #0 ap_CS_fsm = 15'd1;
    #0 ap_enable_reg_pp1_iter0 = 1'b0;
    #0 ap_enable_reg_pp1_iter1 = 1'b0;
  end


  AddRoundKey_Invercud
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  ret_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(ret_address0),
    .ce0(ret_ce0),
    .we0(ret_we0),
    .d0(xor_ln523_reg_1470),
    .q0(ret_q0),
    .address1(ret_address1),
    .ce1(ret_ce1),
    .q1(ret_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_enable_reg_pp1_iter0 <= 1'b0;
    end else
      if((1'b0 == ap_block_pp1_stage0_subdone) & (1'b1 == ap_condition_pp1_exit_iter0_state13) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
        ap_enable_reg_pp1_iter0 <= 1'b0;
      end else if((1'b1 == ap_CS_fsm_state7) & (icmp_ln515_fu_500_p2 == 1'd1)) begin
        ap_enable_reg_pp1_iter0 <= 1'b1;
      end 
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_enable_reg_pp1_iter1 <= 1'b0;
    end else
      if((1'b0 == ap_block_pp1_stage1_subdone) & (1'b1 == ap_CS_fsm_pp1_stage1) | (1'b0 == ap_block_pp1_stage0_subdone) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
        ap_enable_reg_pp1_iter1 <= ap_enable_reg_pp1_iter0;
      end else if((1'b1 == ap_CS_fsm_state7) & (icmp_ln515_fu_500_p2 == 1'd1)) begin
        ap_enable_reg_pp1_iter1 <= 1'b0;
      end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state7) & (icmp_ln515_fu_500_p2 == 1'd1)) begin
      i_1_reg_325 <= 3'd0;
    end else if((icmp_ln526_reg_1475 == 1'd0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      i_1_reg_325 <= i_reg_1479;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln515_fu_500_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      i_assign_reg_314 <= 3'd0;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      i_assign_reg_314 <= i_5_reg_1365;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      j_0_reg_292 <= j_reg_1285;
    end else if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      j_0_reg_292 <= 3'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      j_assign_reg_303 <= 3'd0;
    end else if((1'b1 == ap_CS_fsm_state8) & (icmp_ln516_fu_528_p2 == 1'd1)) begin
      j_assign_reg_303 <= j_1_reg_1345;
    end 
  end

  assign shl_ln_fu_431_p3_temp_6 = shl_ln_fu_431_p3 & 3'd12;
  assign shl_ln_reg_1305_temp_7 = shl_ln_reg_1305 & 3'd3;
  assign shl_ln_fu_431_p3_temp_6_temp_8 = shl_ln_fu_431_p3_temp_6 | shl_ln_reg_1305_temp_7;
  assign zext_ln511_fu_450_p1_temp_9 = zext_ln511_fu_450_p1 & 63'd12;
  assign statemt_addr_17_reg_1316_temp_10 = statemt_addr_17_reg_1316 & 4'd19;
  assign zext_ln511_fu_450_p1_temp_9_temp_11 = zext_ln511_fu_450_p1_temp_9 | statemt_addr_17_reg_1316_temp_10;
  assign zext_ln510_fu_439_p1_temp_12 = zext_ln510_fu_439_p1 & 63'd12;
  assign statemt_addr_reg_1311_temp_13 = statemt_addr_reg_1311 & 4'd19;
  assign zext_ln510_fu_439_p1_temp_12_temp_14 = zext_ln510_fu_439_p1_temp_12 | statemt_addr_reg_1311_temp_13;

  always @(posedge ap_clk) begin
    if((icmp_ln507_fu_386_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      add_ln510_reg_1290 <= add_ln510_fu_402_p2;
      shl_ln_reg_1305 <= shl_ln_fu_431_p3_temp_6_temp_8;
      statemt_addr_17_reg_1316 <= zext_ln511_fu_450_p1_temp_9_temp_11;
      statemt_addr_reg_1311 <= zext_ln510_fu_439_p1_temp_12_temp_14;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      i_5_reg_1365 <= i_5_fu_534_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_enable_reg_pp1_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      i_reg_1479 <= i_fu_1223_p2;
    end 
  end

  assign select_ln457_fu_638_p3_temp_15 = select_ln457_fu_638_p3 >> 1'd7;
  assign select_ln457_fu_638_p3_temp_16 = select_ln457_fu_638_p3_temp_15 & 24'd16777215;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      icmp_ln444_reg_1391 <= icmp_ln444_fu_580_p2;
      select_ln457_reg_1413 <= select_ln457_fu_638_p3;
      statemt_load_20_reg_1407 <= statemt_q1;
      tmp_5_reg_1418 <= select_ln457_fu_638_p3_temp_16;
      trunc_ln445_reg_1396 <= trunc_ln445_fu_586_p1;
      trunc_ln446_reg_1401 <= trunc_ln446_fu_590_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      icmp_ln526_reg_1475 <= icmp_ln526_fu_1217_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      j_1_reg_1345 <= j_1_fu_506_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      j_reg_1285 <= j_fu_392_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3)) begin
      reg_368 <= grp_fu_336_p2;
      reg_373 <= grp_fu_342_p2;
    end 
  end

  assign xor_ln476_fu_941_p2_temp_17 = xor_ln476_fu_941_p2 >> 1'd7;
  assign xor_ln476_fu_941_p2_temp_18 = xor_ln476_fu_941_p2_temp_17 & 24'd16777215;
  assign select_ln486_fu_1001_p3_temp_19 = select_ln486_fu_1001_p3 >> 1'd7;
  assign select_ln486_fu_1001_p3_temp_20 = select_ln486_fu_1001_p3_temp_19 & 24'd16777215;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state10) begin
      select_ln486_reg_1454 <= select_ln486_fu_1001_p3;
      statemt_load_21_reg_1433 <= statemt_q0;
      statemt_load_22_reg_1449 <= statemt_q1;
      tmp_10_reg_1444 <= xor_ln476_fu_941_p2_temp_18;
      tmp_15_reg_1460 <= select_ln486_fu_1001_p3_temp_20;
      xor_ln476_reg_1438 <= xor_ln476_fu_941_p2;
      xor_ln523_3_reg_1465 <= xor_ln523_3_fu_1019_p2;
    end 
  end

  assign shl_ln1_fu_516_p3_temp_21 = shl_ln1_fu_516_p3 & 3'd12;
  assign shl_ln1_reg_1357_temp_22 = shl_ln1_reg_1357 & 3'd3;
  assign shl_ln1_fu_516_p3_temp_21_temp_23 = shl_ln1_fu_516_p3_temp_21 | shl_ln1_reg_1357_temp_22;

  always @(posedge ap_clk) begin
    if((icmp_ln515_fu_500_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      shl_ln1_reg_1357 <= shl_ln1_fu_516_p3_temp_21_temp_23;
      trunc_ln520_reg_1350 <= trunc_ln520_fu_512_p1;
    end 
  end

  assign shl_ln2_fu_1233_p3_temp_24 = shl_ln2_fu_1233_p3 & 3'd12;
  assign shl_ln2_reg_1484_temp_25 = shl_ln2_reg_1484 & 3'd3;
  assign shl_ln2_fu_1233_p3_temp_24_temp_26 = shl_ln2_fu_1233_p3_temp_24 | shl_ln2_reg_1484_temp_25;
  assign zext_ln529_fu_1241_p1_temp_27 = zext_ln529_fu_1241_p1 & 63'd12;
  assign zext_ln529_reg_1490_temp_28 = zext_ln529_reg_1490 & 63'd18446744073709551603;
  assign zext_ln529_fu_1241_p1_temp_27_temp_29 = zext_ln529_fu_1241_p1_temp_27 | zext_ln529_reg_1490_temp_28;
  assign zext_ln530_fu_1252_p1_temp_30 = zext_ln530_fu_1252_p1 & 63'd12;
  assign zext_ln530_reg_1500_temp_31 = zext_ln530_reg_1500 & 63'd18446744073709551603;
  assign zext_ln530_fu_1252_p1_temp_30_temp_32 = zext_ln530_fu_1252_p1_temp_30 | zext_ln530_reg_1500_temp_31;

  always @(posedge ap_clk) begin
    if((icmp_ln526_fu_1217_p2 == 1'd0) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      shl_ln2_reg_1484 <= shl_ln2_fu_1233_p3_temp_24_temp_26;
      zext_ln529_reg_1490 <= zext_ln529_fu_1241_p1_temp_27_temp_29;
      zext_ln530_reg_1500 <= zext_ln530_fu_1252_p1_temp_30_temp_32;
    end 
  end

  assign shl_ln510_1_fu_378_p3_temp_33 = shl_ln510_1_fu_378_p3 & 5'd60;
  assign shl_ln510_1_reg_1277_temp_34 = shl_ln510_1_reg_1277 & 5'd3;
  assign shl_ln510_1_fu_378_p3_temp_33_temp_35 = shl_ln510_1_fu_378_p3_temp_33 | shl_ln510_1_reg_1277_temp_34;

  always @(posedge ap_clk) begin
    if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      shl_ln510_1_reg_1277 <= shl_ln510_1_fu_378_p3_temp_33_temp_35;
    end 
  end

  assign zext_ln512_fu_485_p1_temp_36 = zext_ln512_fu_485_p1 & 63'd12;
  assign statemt_addr_18_reg_1331_temp_37 = statemt_addr_18_reg_1331 & 4'd19;
  assign zext_ln512_fu_485_p1_temp_36_temp_38 = zext_ln512_fu_485_p1_temp_36 | statemt_addr_18_reg_1331_temp_37;
  assign zext_ln513_fu_495_p1_temp_39 = zext_ln513_fu_495_p1 & 63'd12;
  assign statemt_addr_19_reg_1336_temp_40 = statemt_addr_19_reg_1336 & 4'd19;
  assign zext_ln513_fu_495_p1_temp_39_temp_41 = zext_ln513_fu_495_p1_temp_39 | statemt_addr_19_reg_1336_temp_40;

  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_addr_18_reg_1331 <= zext_ln512_fu_485_p1_temp_36_temp_38;
      statemt_addr_19_reg_1336 <= zext_ln513_fu_495_p1_temp_39_temp_41;
    end 
  end

  assign zext_ln443_fu_545_p1_temp_42 = zext_ln443_fu_545_p1 & 4'd15;
  assign zext_ln443_reg_1370_temp_43 = zext_ln443_reg_1370 & 4'd18446744073709551600;
  assign zext_ln443_fu_545_p1_temp_42_temp_44 = zext_ln443_fu_545_p1_temp_42 | zext_ln443_reg_1370_temp_43;

  always @(posedge ap_clk) begin
    if((icmp_ln516_fu_528_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state8)) begin
      trunc_ln456_reg_1380 <= trunc_ln456_fu_550_p1;
      zext_ln443_reg_1370 <= zext_ln443_fu_545_p1_temp_42_temp_44;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      xor_ln523_reg_1470 <= xor_ln523_fu_1211_p2;
    end 
  end

  assign zext_ln531_fu_1262_p1_temp_45 = zext_ln531_fu_1262_p1 & 63'd12;
  assign zext_ln531_reg_1510_temp_46 = zext_ln531_reg_1510 & 63'd18446744073709551603;
  assign zext_ln531_fu_1262_p1_temp_45_temp_47 = zext_ln531_fu_1262_p1_temp_45 | zext_ln531_reg_1510_temp_46;
  assign zext_ln532_fu_1272_p1_temp_48 = zext_ln532_fu_1272_p1 & 63'd12;
  assign zext_ln532_reg_1520_temp_49 = zext_ln532_reg_1520 & 63'd18446744073709551603;
  assign zext_ln532_fu_1272_p1_temp_48_temp_50 = zext_ln532_fu_1272_p1_temp_48 | zext_ln532_reg_1520_temp_49;

  always @(posedge ap_clk) begin
    if((icmp_ln526_reg_1475 == 1'd0) & (1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1)) begin
      zext_ln531_reg_1510 <= zext_ln531_fu_1262_p1_temp_45_temp_47;
      zext_ln532_reg_1520 <= zext_ln532_fu_1272_p1_temp_48_temp_50;
    end 
  end


  always @(*) begin
    if(icmp_ln526_fu_1217_p2 == 1'd1) begin
      ap_condition_pp1_exit_iter0_state13 = 1'b1;
    end else begin
      ap_condition_pp1_exit_iter0_state13 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state16) | (ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((ap_enable_reg_pp1_iter1 == 1'b0) & (ap_enable_reg_pp1_iter0 == 1'b0)) begin
      ap_idle_pp1 = 1'b1;
    end else begin
      ap_idle_pp1 = 1'b0;
    end
  end


  always @(*) begin
    if((icmp_ln526_reg_1475 == 1'd0) & (1'b0 == ap_block_pp1_stage0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
      ap_phi_mux_i_1_phi_fu_329_p4 = i_reg_1479;
    end else begin
      ap_phi_mux_i_1_phi_fu_329_p4 = i_1_reg_325;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_pp1_stage1) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
      ret_address0 = zext_ln532_fu_1272_p1;
    end else if((1'b0 == ap_block_pp1_stage0) & (ap_enable_reg_pp1_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
      ret_address0 = zext_ln529_fu_1241_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      ret_address0 = zext_ln443_reg_1370;
    end else begin
      ret_address0 = 'bx;
    end
  end


  always @(*) begin
      if((1'b0 == ap_block_pp1_stage1) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
        ret_address1 = zext_ln531_fu_1262_p1;
      end else if((1'b0 == ap_block_pp1_stage0) & (1'b1 == ap_CS_fsm_pp1_stage0) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
        ret_address1 = zext_ln530_fu_1252_p1;
      end else if(ap_enable_reg_pp1_iter0 == 1'b1) begin
        ret_address1 = 'bx;
      end else begin
      ret_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state12) | (1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1) | (ap_enable_reg_pp1_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      ret_ce0 = 1'b1;
    end else begin
      ret_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1) | (ap_enable_reg_pp1_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      ret_ce1 = 1'b1;
    end else begin
      ret_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state12) begin
      ret_we0 = 1'b1;
    end else begin
      ret_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_pp1_stage0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
      statemt_address0 = zext_ln531_reg_1510;
    end else if((1'b0 == ap_block_pp1_stage1) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
      statemt_address0 = zext_ln529_reg_1490;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_address0 = zext_ln472_fu_668_p1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = zext_ln443_fu_545_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address0 = statemt_addr_18_reg_1331;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address0 = statemt_addr_reg_1311;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = zext_ln512_fu_485_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address0 = zext_ln510_fu_439_p1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_pp1_stage0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
      statemt_address1 = zext_ln532_reg_1520;
    end else if((1'b0 == ap_block_pp1_stage1) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
      statemt_address1 = zext_ln530_reg_1500;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_address1 = zext_ln485_fu_685_p1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = zext_ln456_fu_567_p1;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address1 = statemt_addr_19_reg_1336;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address1 = statemt_addr_17_reg_1316;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address1 = zext_ln513_fu_495_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address1 = zext_ln511_fu_450_p1;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1) | (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state8) | (1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1) | (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      statemt_ce1 = 1'b1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_pp1_stage0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
      statemt_d0 = ret_q1;
    end else if((1'b0 == ap_block_pp1_stage1) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
      statemt_d0 = ret_q0;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d0 = reg_368;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b0 == ap_block_pp1_stage0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0)) begin
      statemt_d1 = ret_q0;
    end else if((1'b0 == ap_block_pp1_stage1) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1)) begin
      statemt_d1 = ret_q1;
    end else if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5)) begin
      statemt_d1 = reg_373;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5) | (icmp_ln526_reg_1475 == 1'd0) & (1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1) | (icmp_ln526_reg_1475 == 1'd0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state5) | (icmp_ln526_reg_1475 == 1'd0) & (1'b0 == ap_block_pp1_stage1_11001) & (1'b1 == ap_CS_fsm_pp1_stage1) & (ap_enable_reg_pp1_iter0 == 1'b1) | (icmp_ln526_reg_1475 == 1'd0) & (ap_enable_reg_pp1_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp1_stage0) & (1'b0 == ap_block_pp1_stage0_11001)) begin
      statemt_we1 = 1'b1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address0 = zext_ln512_1_fu_464_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address0 = zext_ln510_1_fu_407_p1;
    end else begin
      word_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      word_address1 = zext_ln513_1_fu_475_p1;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      word_address1 = zext_ln511_1_fu_422_p1;
    end else begin
      word_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce0 = 1'b1;
    end else begin
      word_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state3)) begin
      word_ce1 = 1'b1;
    end else begin
      word_ce1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((icmp_ln507_fu_386_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state6: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state7: begin
        if((1'b1 == ap_CS_fsm_state7) & (icmp_ln515_fu_500_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_pp1_stage0;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        if((1'b1 == ap_CS_fsm_state8) & (icmp_ln516_fu_528_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state12: begin
        ap_NS_fsm = ap_ST_fsm_state8;
      end
      ap_ST_fsm_pp1_stage0: begin
        if(~((1'b0 == ap_block_pp1_stage0_subdone) & (ap_enable_reg_pp1_iter0 == 1'b1) & (icmp_ln526_fu_1217_p2 == 1'd1)) & (1'b0 == ap_block_pp1_stage0_subdone)) begin
          ap_NS_fsm = ap_ST_fsm_pp1_stage1;
        end else if((1'b0 == ap_block_pp1_stage0_subdone) & (ap_enable_reg_pp1_iter0 == 1'b1) & (icmp_ln526_fu_1217_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state16;
        end else begin
          ap_NS_fsm = ap_ST_fsm_pp1_stage0;
        end
      end
      ap_ST_fsm_pp1_stage1: begin
        if(1'b0 == ap_block_pp1_stage1_subdone) begin
          ap_NS_fsm = ap_ST_fsm_pp1_stage0;
        end else begin
          ap_NS_fsm = ap_ST_fsm_pp1_stage1;
        end
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state1;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign add_ln443_fu_540_p2 = zext_ln516_fu_524_p1 + shl_ln1_reg_1357;
  assign add_ln456_1_fu_554_p2 = trunc_ln456_fu_550_p1 + 2'd1;
  assign add_ln485_fu_673_p2 = $signed(trunc_ln456_reg_1380) + $signed(2'd3);
  assign add_ln510_fu_402_p2 = zext_ln507_fu_398_p1 + shl_ln510_1_reg_1277;
  assign add_ln511_fu_416_p2 = 8'd120 + zext_ln510_3_fu_412_p1;
  assign add_ln512_fu_458_p2 = 9'd240 + zext_ln510_2_fu_455_p1;
  assign add_ln513_fu_469_p2 = $signed(9'd360) + $signed(zext_ln510_2_fu_455_p1);
  assign tmp_15_reg_1460_temp_51 = tmp_15_reg_1460 << 1'd8;
  assign and_ln10_fu_1108_p3 = tmp_15_reg_1460_temp_51;
  assign tmp_16_fu_1153_p4_temp_52 = tmp_16_fu_1153_p4 << 1'd8;
  assign and_ln11_fu_1163_p3 = tmp_16_fu_1153_p4_temp_52;
  assign tmp_8_fu_715_p4_temp_53 = tmp_8_fu_715_p4 << 1'd8;
  assign and_ln1_fu_725_p3 = tmp_8_fu_715_p4_temp_53;
  assign tmp_s_fu_772_p4_temp_54 = tmp_s_fu_772_p4 << 1'd8;
  assign and_ln2_fu_782_p3 = tmp_s_fu_772_p4_temp_54;
  assign grp_fu_358_p4_temp_55 = grp_fu_358_p4 << 1'd8;
  assign and_ln3_fu_594_p3 = grp_fu_358_p4_temp_55;
  assign tmp_5_reg_1418_temp_56 = tmp_5_reg_1418 << 1'd8;
  assign and_ln4_fu_813_p3 = tmp_5_reg_1418_temp_56;
  assign tmp_7_fu_859_p4_temp_57 = tmp_7_fu_859_p4 << 1'd8;
  assign and_ln5_fu_869_p3 = tmp_7_fu_859_p4_temp_57;
  assign grp_fu_348_p4_temp_58 = grp_fu_348_p4 << 1'd8;
  assign and_ln6_fu_897_p3 = grp_fu_348_p4_temp_58;
  assign tmp_10_reg_1444_temp_59 = tmp_10_reg_1444 << 1'd8;
  assign and_ln7_fu_1025_p3 = tmp_10_reg_1444_temp_59;
  assign tmp_11_fu_1070_p4_temp_60 = tmp_11_fu_1070_p4 << 1'd8;
  assign and_ln8_fu_1080_p3 = tmp_11_fu_1070_p4_temp_60;
  assign grp_fu_358_p4_temp_61 = grp_fu_358_p4 << 1'd8;
  assign and_ln9_fu_957_p3 = grp_fu_358_p4_temp_61;
  assign grp_fu_348_p4_temp_62 = grp_fu_348_p4 << 1'd8;
  assign and_ln_fu_572_p3 = grp_fu_348_p4_temp_62;
  assign ap_CS_fsm_pp1_stage0 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_pp1_stage1 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign ap_block_pp1_stage0 = ~(1'b1 == 1'b1);
  assign ap_block_pp1_stage0_11001 = ~(1'b1 == 1'b1);
  assign ap_block_pp1_stage0_subdone = ~(1'b1 == 1'b1);
  assign ap_block_pp1_stage1 = ~(1'b1 == 1'b1);
  assign ap_block_pp1_stage1_11001 = ~(1'b1 == 1'b1);
  assign ap_block_pp1_stage1_subdone = ~(1'b1 == 1'b1);
  assign ap_block_state13_pp1_stage0_iter0 = ~(1'b1 == 1'b1);
  assign ap_block_state14_pp1_stage1_iter0 = ~(1'b1 == 1'b1);
  assign ap_block_state15_pp1_stage0_iter1 = ~(1'b1 == 1'b1);
  assign ap_enable_pp1 = ap_idle_pp1 ^ 1'b1;
  assign grp_fu_336_p2 = word_q0 ^ statemt_q0;
  assign grp_fu_342_p2 = word_q1 ^ statemt_q1;
  assign statemt_q0_temp_63 = statemt_q0 >> 1'd7;
  assign statemt_q0_temp_64 = statemt_q0_temp_63 & 24'd16777215;
  assign grp_fu_348_p4 = statemt_q0_temp_64;
  assign statemt_q1_temp_65 = statemt_q1 >> 1'd7;
  assign statemt_q1_temp_66 = statemt_q1_temp_65 & 24'd16777215;
  assign grp_fu_358_p4 = statemt_q1_temp_66;
  assign i_5_fu_534_p2 = i_assign_reg_314 + 3'd1;
  assign i_fu_1223_p2 = ap_phi_mux_i_1_phi_fu_329_p4 + 3'd1;
  assign icmp_ln444_fu_580_p2 = (and_ln_fu_572_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln448_fu_733_p2 = (and_ln1_fu_725_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln452_fu_790_p2 = (and_ln2_fu_782_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln457_fu_602_p2 = (and_ln3_fu_594_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln460_fu_820_p2 = (and_ln4_fu_813_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln464_fu_877_p2 = (and_ln5_fu_869_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln473_fu_905_p2 = (and_ln6_fu_897_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln477_fu_1032_p2 = (and_ln7_fu_1025_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln480_fu_1088_p2 = (and_ln8_fu_1080_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln486_fu_965_p2 = (and_ln9_fu_957_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln489_fu_1115_p2 = (and_ln10_fu_1108_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln492_fu_1171_p2 = (and_ln11_fu_1163_p3 == 32'd256)? 1'b1 : 1'b0;
  assign icmp_ln507_fu_386_p2 = (j_0_reg_292 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln515_fu_500_p2 = (j_assign_reg_303 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln516_fu_528_p2 = (i_assign_reg_314 == 3'd4)? 1'b1 : 1'b0;
  assign icmp_ln526_fu_1217_p2 = (ap_phi_mux_i_1_phi_fu_329_p4 == 3'd4)? 1'b1 : 1'b0;
  assign j_1_fu_506_p2 = j_assign_reg_303 + 3'd1;
  assign j_fu_392_p2 = j_0_reg_292 + 3'd1;
  assign trunc_ln520_reg_1350_temp_67 = trunc_ln520_reg_1350 << 1'd2;
  assign trunc_ln520_reg_1350_temp_68 = trunc_ln520_reg_1350_temp_67 | xor_ln472_fu_656_p2;
  assign or_ln1_fu_661_p3 = trunc_ln520_reg_1350_temp_68;
  assign trunc_ln520_reg_1350_temp_69 = trunc_ln520_reg_1350 << 1'd2;
  assign trunc_ln520_reg_1350_temp_70 = trunc_ln520_reg_1350_temp_69 | add_ln485_fu_673_p2;
  assign or_ln2_fu_678_p3 = trunc_ln520_reg_1350_temp_70;
  assign or_ln511_fu_444_p2 = shl_ln_fu_431_p3 | 4'd1;
  assign or_ln512_fu_480_p2 = shl_ln_reg_1305 | 4'd2;
  assign or_ln513_fu_490_p2 = shl_ln_reg_1305 | 4'd3;
  assign or_ln530_fu_1246_p2 = shl_ln2_fu_1233_p3 | 4'd1;
  assign or_ln531_fu_1257_p2 = shl_ln2_reg_1484 | 4'd2;
  assign or_ln532_fu_1267_p2 = shl_ln2_reg_1484 | 4'd3;
  assign trunc_ln520_reg_1350_temp_71 = trunc_ln520_reg_1350 << 1'd2;
  assign trunc_ln520_reg_1350_temp_72 = trunc_ln520_reg_1350_temp_71 | add_ln456_1_fu_554_p2;
  assign or_ln_fu_560_p3 = trunc_ln520_reg_1350_temp_72;
  assign icmp_ln444_reg_1391_temp_73 = icmp_ln444_reg_1391 & 30'd1;
  assign select_ln444_fu_703_p3 = (icmp_ln444_reg_1391_temp_73 === 1'b1)? xor_ln444_fu_697_p2 : trunc_ln_fu_690_p3;
  assign icmp_ln448_fu_733_p2_temp_74 = icmp_ln448_fu_733_p2 & 30'd1;
  assign select_ln448_fu_751_p3 = (icmp_ln448_fu_733_p2_temp_74 === 1'b1)? xor_ln448_fu_745_p2 : shl_ln449_fu_739_p2;
  assign icmp_ln452_fu_790_p2_temp_75 = icmp_ln452_fu_790_p2 & 31'd1;
  assign select_ln452_fu_802_p3 = (icmp_ln452_fu_790_p2_temp_75 === 1'b1)? xor_ln453_fu_796_p2 : x_assign_2_fu_764_p3;
  assign icmp_ln457_fu_602_p2_temp_76 = icmp_ln457_fu_602_p2 & 30'd1;
  assign select_ln457_fu_638_p3 = (icmp_ln457_fu_602_p2_temp_76 === 1'b1)? xor_ln459_fu_620_p2 : tmp_4_fu_630_p3;
  assign icmp_ln460_fu_820_p2_temp_77 = icmp_ln460_fu_820_p2 & 30'd1;
  assign select_ln460_fu_837_p3 = (icmp_ln460_fu_820_p2_temp_77 === 1'b1)? xor_ln460_fu_831_p2 : shl_ln461_fu_826_p2;
  assign icmp_ln464_fu_877_p2_temp_78 = icmp_ln464_fu_877_p2 & 31'd1;
  assign select_ln464_fu_889_p3 = (icmp_ln464_fu_877_p2_temp_78 === 1'b1)? xor_ln465_fu_883_p2 : x_assign_9_fu_851_p3;
  assign icmp_ln473_fu_905_p2_temp_79 = icmp_ln473_fu_905_p2 & 30'd1;
  assign select_ln473_fu_929_p3 = (icmp_ln473_fu_905_p2_temp_79 === 1'b1)? xor_ln473_fu_923_p2 : trunc_ln6_fu_915_p3;
  assign icmp_ln477_fu_1032_p2_temp_80 = icmp_ln477_fu_1032_p2 & 30'd1;
  assign select_ln477_fu_1054_p3 = (icmp_ln477_fu_1032_p2_temp_80 === 1'b1)? xor_ln479_fu_1043_p2 : shl_ln479_fu_1049_p2;
  assign icmp_ln480_fu_1088_p2_temp_81 = icmp_ln480_fu_1088_p2 & 31'd1;
  assign select_ln480_fu_1100_p3 = (icmp_ln480_fu_1088_p2_temp_81 === 1'b1)? xor_ln481_fu_1094_p2 : x_assign_1_fu_1062_p3;
  assign icmp_ln486_fu_965_p2_temp_82 = icmp_ln486_fu_965_p2 & 30'd1;
  assign select_ln486_fu_1001_p3 = (icmp_ln486_fu_965_p2_temp_82 === 1'b1)? xor_ln488_fu_983_p2 : tmp_14_fu_993_p3;
  assign icmp_ln489_fu_1115_p2_temp_83 = icmp_ln489_fu_1115_p2 & 30'd1;
  assign select_ln489_fu_1137_p3 = (icmp_ln489_fu_1115_p2_temp_83 === 1'b1)? xor_ln491_fu_1126_p2 : shl_ln491_fu_1132_p2;
  assign icmp_ln492_fu_1171_p2_temp_84 = icmp_ln492_fu_1171_p2 & 31'd1;
  assign select_ln492_fu_1183_p3 = (icmp_ln492_fu_1171_p2_temp_84 === 1'b1)? xor_ln493_fu_1177_p2 : x_assign_6_fu_1145_p3;
  assign trunc_ln520_fu_512_p1_temp_85 = trunc_ln520_fu_512_p1 << 1'd2;
  assign shl_ln1_fu_516_p3 = trunc_ln520_fu_512_p1_temp_85;
  assign trunc_ln529_fu_1229_p1_temp_86 = trunc_ln529_fu_1229_p1 << 1'd2;
  assign shl_ln2_fu_1233_p3 = trunc_ln529_fu_1229_p1_temp_86;
  assign shl_ln449_fu_739_p2 = xor_ln447_fu_710_p2 << 31'd1;
  assign shl_ln461_fu_826_p2 = select_ln457_reg_1413 << 31'd1;
  assign shl_ln478_fu_1038_p2 = xor_ln476_reg_1438 << 31'd1;
  assign shl_ln479_fu_1049_p2 = xor_ln476_reg_1438 << 31'd1;
  assign shl_ln490_fu_1121_p2 = select_ln486_reg_1454 << 31'd1;
  assign shl_ln491_fu_1132_p2 = select_ln486_reg_1454 << 31'd1;
  assign n_temp_87 = n << 1'd2;
  assign shl_ln510_1_fu_378_p3 = n_temp_87;
  assign trunc_ln510_fu_427_p1_temp_88 = trunc_ln510_fu_427_p1 << 1'd2;
  assign shl_ln_fu_431_p3 = trunc_ln510_fu_427_p1_temp_88;
  assign select_ln477_fu_1054_p3_temp_89 = select_ln477_fu_1054_p3 >> 1'd7;
  assign select_ln477_fu_1054_p3_temp_90 = select_ln477_fu_1054_p3_temp_89 & 24'd16777215;
  assign tmp_11_fu_1070_p4 = select_ln477_fu_1054_p3_temp_90;
  assign trunc_ln487_fu_971_p1_temp_91 = trunc_ln487_fu_971_p1 << 1'd1;
  assign tmp_13_fu_975_p3 = trunc_ln487_fu_971_p1_temp_91;
  assign trunc_ln488_fu_989_p1_temp_92 = trunc_ln488_fu_989_p1 << 1'd1;
  assign tmp_14_fu_993_p3 = trunc_ln488_fu_989_p1_temp_92;
  assign select_ln489_fu_1137_p3_temp_93 = select_ln489_fu_1137_p3 >> 1'd7;
  assign select_ln489_fu_1137_p3_temp_94 = select_ln489_fu_1137_p3_temp_93 & 24'd16777215;
  assign tmp_16_fu_1153_p4 = select_ln489_fu_1137_p3_temp_94;
  assign trunc_ln458_fu_608_p1_temp_95 = trunc_ln458_fu_608_p1 << 1'd1;
  assign tmp_3_fu_612_p3 = trunc_ln458_fu_608_p1_temp_95;
  assign trunc_ln459_fu_626_p1_temp_96 = trunc_ln459_fu_626_p1 << 1'd1;
  assign tmp_4_fu_630_p3 = trunc_ln459_fu_626_p1_temp_96;
  assign xor_ln463_fu_845_p2_temp_97 = xor_ln463_fu_845_p2 >> 1'd7;
  assign xor_ln463_fu_845_p2_temp_98 = xor_ln463_fu_845_p2_temp_97 & 24'd16777215;
  assign tmp_7_fu_859_p4 = xor_ln463_fu_845_p2_temp_98;
  assign xor_ln447_fu_710_p2_temp_99 = xor_ln447_fu_710_p2 >> 1'd7;
  assign xor_ln447_fu_710_p2_temp_100 = xor_ln447_fu_710_p2_temp_99 & 24'd16777215;
  assign tmp_8_fu_715_p4 = xor_ln447_fu_710_p2_temp_100;
  assign xor_ln451_fu_759_p2_temp_101 = xor_ln451_fu_759_p2 >> 1'd7;
  assign xor_ln451_fu_759_p2_temp_102 = xor_ln451_fu_759_p2_temp_101 & 24'd16777215;
  assign tmp_s_fu_772_p4 = xor_ln451_fu_759_p2_temp_102;
  assign trunc_ln445_fu_586_p1 = (statemt_q0 & 30'd1073741823);
  assign trunc_ln446_fu_590_p1 = (statemt_q0 & 31'd2147483647);
  assign trunc_ln456_1_fu_810_p1 = (statemt_load_20_reg_1407 & 31'd2147483647);
  assign trunc_ln456_fu_550_p1 = (i_assign_reg_314 & 2'd3);
  assign trunc_ln458_fu_608_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln459_fu_626_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln474_fu_911_p1 = (statemt_q0 & 30'd1073741823);
  assign trunc_ln475_fu_937_p1 = (statemt_q0 & 31'd2147483647);
  assign trunc_ln487_fu_971_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln488_fu_989_p1 = (statemt_q1 & 30'd1073741823);
  assign trunc_ln510_fu_427_p1 = (j_0_reg_292 & 2'd3);
  assign trunc_ln520_fu_512_p1 = (j_assign_reg_303 & 2'd3);
  assign trunc_ln529_fu_1229_p1 = (ap_phi_mux_i_1_phi_fu_329_p4 & 2'd3);
  assign trunc_ln474_fu_911_p1_temp_103 = trunc_ln474_fu_911_p1 << 1'd1;
  assign trunc_ln6_fu_915_p3 = trunc_ln474_fu_911_p1_temp_103;
  assign trunc_ln445_reg_1396_temp_104 = trunc_ln445_reg_1396 << 1'd1;
  assign trunc_ln_fu_690_p3 = trunc_ln445_reg_1396_temp_104;
  assign select_ln477_fu_1054_p3_temp_105 = select_ln477_fu_1054_p3 << 1'd1;
  assign x_assign_1_fu_1062_p3 = select_ln477_fu_1054_p3_temp_105;
  assign xor_ln451_fu_759_p2_temp_106 = xor_ln451_fu_759_p2 << 1'd1;
  assign x_assign_2_fu_764_p3 = xor_ln451_fu_759_p2_temp_106;
  assign select_ln489_fu_1137_p3_temp_107 = select_ln489_fu_1137_p3 << 1'd1;
  assign x_assign_6_fu_1145_p3 = select_ln489_fu_1137_p3_temp_107;
  assign xor_ln463_fu_845_p2_temp_108 = xor_ln463_fu_845_p2 << 1'd1;
  assign x_assign_9_fu_851_p3 = xor_ln463_fu_845_p2_temp_108;
  assign xor_ln444_fu_697_p2 = trunc_ln_fu_690_p3 ^ 31'd283;
  assign xor_ln447_fu_710_p2 = trunc_ln446_reg_1401 ^ select_ln444_fu_703_p3;
  assign xor_ln448_fu_745_p2 = shl_ln449_fu_739_p2 ^ 31'd283;
  assign xor_ln451_fu_759_p2 = trunc_ln446_reg_1401 ^ select_ln448_fu_751_p3;
  assign xor_ln453_fu_796_p2 = x_assign_2_fu_764_p3 ^ 32'd283;
  assign xor_ln459_fu_620_p2 = tmp_3_fu_612_p3 ^ 31'd283;
  assign xor_ln460_fu_831_p2 = shl_ln461_fu_826_p2 ^ 31'd283;
  assign xor_ln463_fu_845_p2 = trunc_ln456_1_fu_810_p1 ^ select_ln460_fu_837_p3;
  assign xor_ln465_fu_883_p2 = x_assign_9_fu_851_p3 ^ 32'd283;
  assign xor_ln472_fu_656_p2 = trunc_ln456_reg_1380 ^ 2'd2;
  assign xor_ln473_fu_923_p2 = trunc_ln6_fu_915_p3 ^ 31'd283;
  assign xor_ln476_fu_941_p2 = trunc_ln475_fu_937_p1 ^ select_ln473_fu_929_p3;
  assign xor_ln479_fu_1043_p2 = shl_ln478_fu_1038_p2 ^ 31'd283;
  assign xor_ln481_fu_1094_p2 = x_assign_1_fu_1062_p3 ^ 32'd283;
  assign xor_ln488_fu_983_p2 = tmp_13_fu_975_p3 ^ 31'd283;
  assign xor_ln491_fu_1126_p2 = shl_ln490_fu_1121_p2 ^ 31'd283;
  assign xor_ln493_fu_1177_p2 = x_assign_6_fu_1145_p3 ^ 32'd283;
  assign xor_ln523_1_fu_1191_p2 = statemt_load_22_reg_1449 ^ statemt_load_21_reg_1433;
  assign xor_ln523_2_fu_1195_p2 = xor_ln523_1_fu_1191_p2 ^ statemt_load_20_reg_1407;
  assign xor_ln523_3_fu_1019_p2 = select_ln464_fu_889_p3 ^ select_ln452_fu_802_p3;
  assign xor_ln523_4_fu_1200_p2 = select_ln492_fu_1183_p3 ^ select_ln480_fu_1100_p3;
  assign xor_ln523_5_fu_1206_p2 = xor_ln523_4_fu_1200_p2 ^ xor_ln523_3_reg_1465;
  assign xor_ln523_fu_1211_p2 = xor_ln523_5_fu_1206_p2 ^ xor_ln523_2_fu_1195_p2;
  assign zext_ln443_fu_545_p1 = add_ln443_fu_540_p2;
  assign zext_ln456_fu_567_p1 = or_ln_fu_560_p3;
  assign zext_ln472_fu_668_p1 = or_ln1_fu_661_p3;
  assign zext_ln485_fu_685_p1 = or_ln2_fu_678_p3;
  assign zext_ln507_fu_398_p1 = j_0_reg_292;
  assign zext_ln510_1_fu_407_p1 = add_ln510_fu_402_p2;
  assign zext_ln510_2_fu_455_p1 = add_ln510_reg_1290;
  assign zext_ln510_3_fu_412_p1 = add_ln510_fu_402_p2;
  assign zext_ln510_fu_439_p1 = shl_ln_fu_431_p3;
  assign zext_ln511_1_fu_422_p1 = add_ln511_fu_416_p2;
  assign zext_ln511_fu_450_p1 = or_ln511_fu_444_p2;
  assign zext_ln512_1_fu_464_p1 = add_ln512_fu_458_p2;
  assign zext_ln512_fu_485_p1 = or_ln512_fu_480_p2;
  assign zext_ln513_1_fu_475_p1 = add_ln513_fu_469_p2;
  assign zext_ln513_fu_495_p1 = or_ln513_fu_490_p2;
  assign zext_ln516_fu_524_p1 = i_assign_reg_314;
  assign zext_ln529_fu_1241_p1 = shl_ln2_fu_1233_p3;
  assign zext_ln530_fu_1252_p1 = or_ln530_fu_1246_p2;
  assign zext_ln531_fu_1262_p1 = or_ln531_fu_1257_p2;
  assign zext_ln532_fu_1272_p1 = or_ln532_fu_1267_p2;

  always @(posedge ap_clk) begin
    shl_ln510_1_reg_1277 <= shl_ln510_1_reg_1277 & 1'd60;
    shl_ln_reg_1305 <= shl_ln_reg_1305 & 1'd12;
    statemt_addr_reg_1311 <= statemt_addr_reg_1311 & 1'd28;
    statemt_addr_reg_1311 <= statemt_addr_reg_1311 & 4'd15;
    statemt_addr_17_reg_1316 <= statemt_addr_17_reg_1316 & 1'd29;
    statemt_addr_17_reg_1316 <= statemt_addr_17_reg_1316 & 4'd15;
    statemt_addr_18_reg_1331 <= statemt_addr_18_reg_1331 & 1'd30;
    statemt_addr_18_reg_1331 <= statemt_addr_18_reg_1331 & 4'd15;
    statemt_addr_19_reg_1336 <= statemt_addr_19_reg_1336 & 1'd31;
    statemt_addr_19_reg_1336 <= statemt_addr_19_reg_1336 & 4'd15;
    shl_ln1_reg_1357 <= shl_ln1_reg_1357 & 1'd12;
    zext_ln443_reg_1370 <= zext_ln443_reg_1370 & 63'd15;
    shl_ln2_reg_1484 <= shl_ln2_reg_1484 & 1'd12;
    zext_ln529_reg_1490 <= zext_ln529_reg_1490 & 1'd18446744073709551612;
    zext_ln529_reg_1490 <= zext_ln529_reg_1490 & 63'd15;
    zext_ln530_reg_1500 <= zext_ln530_reg_1500 & 1'd18446744073709551613;
    zext_ln530_reg_1500 <= zext_ln530_reg_1500 & 63'd15;
    zext_ln531_reg_1510 <= zext_ln531_reg_1510 & 1'd18446744073709551614;
    zext_ln531_reg_1510 <= zext_ln531_reg_1510 & 63'd15;
    zext_ln532_reg_1520 <= zext_ln532_reg_1520 & 1'd18446744073709551615;
    zext_ln532_reg_1520 <= zext_ln532_reg_1520 & 63'd15;
  end


endmodule

