
module aes_decrypt_call
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt1_address0,
  statemt1_ce0,
  statemt1_we0,
  statemt1_d0,
  statemt1_q0,
  statemt1_address1,
  statemt1_ce1,
  statemt1_we1,
  statemt1_d1
);

  parameter ap_ST_fsm_state1 = 28'd1;
  parameter ap_ST_fsm_state2 = 28'd2;
  parameter ap_ST_fsm_state3 = 28'd4;
  parameter ap_ST_fsm_state4 = 28'd8;
  parameter ap_ST_fsm_state5 = 28'd16;
  parameter ap_ST_fsm_state6 = 28'd32;
  parameter ap_ST_fsm_state7 = 28'd64;
  parameter ap_ST_fsm_state8 = 28'd128;
  parameter ap_ST_fsm_state9 = 28'd256;
  parameter ap_ST_fsm_state10 = 28'd512;
  parameter ap_ST_fsm_state11 = 28'd1024;
  parameter ap_ST_fsm_state12 = 28'd2048;
  parameter ap_ST_fsm_state13 = 28'd4096;
  parameter ap_ST_fsm_state14 = 28'd8192;
  parameter ap_ST_fsm_state15 = 28'd16384;
  parameter ap_ST_fsm_state16 = 28'd32768;
  parameter ap_ST_fsm_state17 = 28'd65536;
  parameter ap_ST_fsm_state18 = 28'd131072;
  parameter ap_ST_fsm_state19 = 28'd262144;
  parameter ap_ST_fsm_state20 = 28'd524288;
  parameter ap_ST_fsm_state21 = 28'd1048576;
  parameter ap_ST_fsm_state22 = 28'd2097152;
  parameter ap_ST_fsm_state23 = 28'd4194304;
  parameter ap_ST_fsm_state24 = 28'd8388608;
  parameter ap_ST_fsm_state25 = 28'd16777216;
  parameter ap_ST_fsm_state26 = 28'd33554432;
  parameter ap_ST_fsm_state27 = 28'd67108864;
  parameter ap_ST_fsm_state28 = 28'd134217728;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt1_address0;
  output statemt1_ce0;
  output statemt1_we0;
  output [31:0] statemt1_d0;
  input [31:0] statemt1_q0;
  output [4:0] statemt1_address1;
  output statemt1_ce1;
  output statemt1_we1;
  output [31:0] statemt1_d1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt1_address0;
  reg statemt1_ce0;
  reg statemt1_we0;
  reg [4:0] statemt1_address1;
  reg statemt1_ce1;
  reg statemt1_we1;
  reg [27:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  wire [31:0] statemt_q0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  wire [31:0] statemt_q1;
  reg [8:0] word_address0;
  reg word_ce0;
  wire [31:0] word_q0;
  reg [8:0] word_address1;
  reg word_ce1;
  wire [31:0] word_q1;
  wire [5:0] i_fu_583_p2;
  reg [5:0] i_reg_609;
  wire ap_CS_fsm_state2;
  wire [63:0] zext_ln12_fu_589_p1;
  reg [63:0] zext_ln12_reg_614;
  wire [0:0] icmp_ln11_fu_577_p2;
  wire [3:0] i_2_fu_600_p2;
  reg [3:0] i_2_reg_627;
  wire ap_CS_fsm_state7;
  wire [0:0] icmp_ln21_fu_594_p2;
  wire grp_AddRoundKey_InversMi_fu_548_ap_start;
  wire grp_AddRoundKey_InversMi_fu_548_ap_done;
  wire grp_AddRoundKey_InversMi_fu_548_ap_idle;
  wire grp_AddRoundKey_InversMi_fu_548_ap_ready;
  wire [4:0] grp_AddRoundKey_InversMi_fu_548_statemt_address0;
  wire grp_AddRoundKey_InversMi_fu_548_statemt_ce0;
  wire grp_AddRoundKey_InversMi_fu_548_statemt_we0;
  wire [31:0] grp_AddRoundKey_InversMi_fu_548_statemt_d0;
  wire [4:0] grp_AddRoundKey_InversMi_fu_548_statemt_address1;
  wire grp_AddRoundKey_InversMi_fu_548_statemt_ce1;
  wire grp_AddRoundKey_InversMi_fu_548_statemt_we1;
  wire [31:0] grp_AddRoundKey_InversMi_fu_548_statemt_d1;
  wire [8:0] grp_AddRoundKey_InversMi_fu_548_word_address0;
  wire grp_AddRoundKey_InversMi_fu_548_word_ce0;
  wire [8:0] grp_AddRoundKey_InversMi_fu_548_word_address1;
  wire grp_AddRoundKey_InversMi_fu_548_word_ce1;
  wire grp_AddRoundKey_fu_558_ap_start;
  wire grp_AddRoundKey_fu_558_ap_done;
  wire grp_AddRoundKey_fu_558_ap_idle;
  wire grp_AddRoundKey_fu_558_ap_ready;
  wire [4:0] grp_AddRoundKey_fu_558_statemt_address0;
  wire grp_AddRoundKey_fu_558_statemt_ce0;
  wire grp_AddRoundKey_fu_558_statemt_we0;
  wire [31:0] grp_AddRoundKey_fu_558_statemt_d0;
  wire [4:0] grp_AddRoundKey_fu_558_statemt_address1;
  wire grp_AddRoundKey_fu_558_statemt_ce1;
  wire grp_AddRoundKey_fu_558_statemt_we1;
  wire [31:0] grp_AddRoundKey_fu_558_statemt_d1;
  reg [4:0] grp_AddRoundKey_fu_558_n;
  wire [8:0] grp_AddRoundKey_fu_558_word_address0;
  wire grp_AddRoundKey_fu_558_word_ce0;
  wire [8:0] grp_AddRoundKey_fu_558_word_address1;
  wire grp_AddRoundKey_fu_558_word_ce1;
  wire grp_InversShiftRow_ByteS_fu_569_ap_start;
  wire grp_InversShiftRow_ByteS_fu_569_ap_done;
  wire grp_InversShiftRow_ByteS_fu_569_ap_idle;
  wire grp_InversShiftRow_ByteS_fu_569_ap_ready;
  wire [4:0] grp_InversShiftRow_ByteS_fu_569_statemt_address0;
  wire grp_InversShiftRow_ByteS_fu_569_statemt_ce0;
  wire grp_InversShiftRow_ByteS_fu_569_statemt_we0;
  wire [31:0] grp_InversShiftRow_ByteS_fu_569_statemt_d0;
  wire [4:0] grp_InversShiftRow_ByteS_fu_569_statemt_address1;
  wire grp_InversShiftRow_ByteS_fu_569_statemt_ce1;
  wire grp_InversShiftRow_ByteS_fu_569_statemt_we1;
  wire [31:0] grp_InversShiftRow_ByteS_fu_569_statemt_d1;
  reg [5:0] i_0_reg_525;
  wire ap_CS_fsm_state3;
  reg [3:0] i_1_reg_536;
  wire ap_CS_fsm_state6;
  wire ap_CS_fsm_state10;
  reg grp_AddRoundKey_InversMi_fu_548_ap_start_reg;
  wire ap_CS_fsm_state8;
  reg grp_AddRoundKey_fu_558_ap_start_reg;
  wire ap_CS_fsm_state4;
  wire ap_CS_fsm_state11;
  reg grp_InversShiftRow_ByteS_fu_569_ap_start_reg;
  wire ap_CS_fsm_state5;
  wire ap_CS_fsm_state9;
  wire ap_CS_fsm_state13;
  wire ap_CS_fsm_state14;
  wire ap_CS_fsm_state15;
  wire ap_CS_fsm_state16;
  wire ap_CS_fsm_state17;
  wire ap_CS_fsm_state18;
  wire ap_CS_fsm_state19;
  wire ap_CS_fsm_state20;
  wire ap_CS_fsm_state21;
  wire ap_CS_fsm_state22;
  wire ap_CS_fsm_state23;
  wire ap_CS_fsm_state24;
  wire ap_CS_fsm_state25;
  wire ap_CS_fsm_state26;
  wire ap_CS_fsm_state27;
  wire ap_CS_fsm_state28;
  wire ap_CS_fsm_state12;
  reg [27:0] ap_NS_fsm;

  initial begin
    #0 ap_CS_fsm = 28'd1;
    #0 grp_AddRoundKey_InversMi_fu_548_ap_start_reg = 1'b0;
    #0 grp_AddRoundKey_fu_558_ap_start_reg = 1'b0;
    #0 grp_InversShiftRow_ByteS_fu_569_ap_start_reg = 1'b0;
  end


  aes_decrypt_call_dEe
  #(
    .DataWidth(32),
    .AddressRange(32),
    .AddressWidth(5)
  )
  statemt_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(statemt_address0),
    .ce0(statemt_ce0),
    .we0(statemt_we0),
    .d0(statemt_d0),
    .q0(statemt_q0),
    .address1(statemt_address1),
    .ce1(statemt_ce1),
    .we1(statemt_we1),
    .d1(statemt_d1),
    .q1(statemt_q1)
  );


  aes_decrypt_call_eOg
  #(
    .DataWidth(32),
    .AddressRange(480),
    .AddressWidth(9)
  )
  word_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(word_address0),
    .ce0(word_ce0),
    .q0(word_q0),
    .address1(word_address1),
    .ce1(word_ce1),
    .q1(word_q1)
  );


  AddRoundKey_InversMi
  grp_AddRoundKey_InversMi_fu_548
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_AddRoundKey_InversMi_fu_548_ap_start),
    .ap_done(grp_AddRoundKey_InversMi_fu_548_ap_done),
    .ap_idle(grp_AddRoundKey_InversMi_fu_548_ap_idle),
    .ap_ready(grp_AddRoundKey_InversMi_fu_548_ap_ready),
    .statemt_address0(grp_AddRoundKey_InversMi_fu_548_statemt_address0),
    .statemt_ce0(grp_AddRoundKey_InversMi_fu_548_statemt_ce0),
    .statemt_we0(grp_AddRoundKey_InversMi_fu_548_statemt_we0),
    .statemt_d0(grp_AddRoundKey_InversMi_fu_548_statemt_d0),
    .statemt_q0(statemt_q0),
    .statemt_address1(grp_AddRoundKey_InversMi_fu_548_statemt_address1),
    .statemt_ce1(grp_AddRoundKey_InversMi_fu_548_statemt_ce1),
    .statemt_we1(grp_AddRoundKey_InversMi_fu_548_statemt_we1),
    .statemt_d1(grp_AddRoundKey_InversMi_fu_548_statemt_d1),
    .statemt_q1(statemt_q1),
    .n(i_1_reg_536),
    .word_address0(grp_AddRoundKey_InversMi_fu_548_word_address0),
    .word_ce0(grp_AddRoundKey_InversMi_fu_548_word_ce0),
    .word_q0(word_q0),
    .word_address1(grp_AddRoundKey_InversMi_fu_548_word_address1),
    .word_ce1(grp_AddRoundKey_InversMi_fu_548_word_ce1),
    .word_q1(word_q1)
  );


  AddRoundKey
  grp_AddRoundKey_fu_558
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_AddRoundKey_fu_558_ap_start),
    .ap_done(grp_AddRoundKey_fu_558_ap_done),
    .ap_idle(grp_AddRoundKey_fu_558_ap_idle),
    .ap_ready(grp_AddRoundKey_fu_558_ap_ready),
    .statemt_address0(grp_AddRoundKey_fu_558_statemt_address0),
    .statemt_ce0(grp_AddRoundKey_fu_558_statemt_ce0),
    .statemt_we0(grp_AddRoundKey_fu_558_statemt_we0),
    .statemt_d0(grp_AddRoundKey_fu_558_statemt_d0),
    .statemt_q0(statemt_q0),
    .statemt_address1(grp_AddRoundKey_fu_558_statemt_address1),
    .statemt_ce1(grp_AddRoundKey_fu_558_statemt_ce1),
    .statemt_we1(grp_AddRoundKey_fu_558_statemt_we1),
    .statemt_d1(grp_AddRoundKey_fu_558_statemt_d1),
    .statemt_q1(statemt_q1),
    .n(grp_AddRoundKey_fu_558_n),
    .word_address0(grp_AddRoundKey_fu_558_word_address0),
    .word_ce0(grp_AddRoundKey_fu_558_word_ce0),
    .word_q0(word_q0),
    .word_address1(grp_AddRoundKey_fu_558_word_address1),
    .word_ce1(grp_AddRoundKey_fu_558_word_ce1),
    .word_q1(word_q1)
  );


  InversShiftRow_ByteS
  grp_InversShiftRow_ByteS_fu_569
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_InversShiftRow_ByteS_fu_569_ap_start),
    .ap_done(grp_InversShiftRow_ByteS_fu_569_ap_done),
    .ap_idle(grp_InversShiftRow_ByteS_fu_569_ap_idle),
    .ap_ready(grp_InversShiftRow_ByteS_fu_569_ap_ready),
    .statemt_address0(grp_InversShiftRow_ByteS_fu_569_statemt_address0),
    .statemt_ce0(grp_InversShiftRow_ByteS_fu_569_statemt_ce0),
    .statemt_we0(grp_InversShiftRow_ByteS_fu_569_statemt_we0),
    .statemt_d0(grp_InversShiftRow_ByteS_fu_569_statemt_d0),
    .statemt_q0(statemt_q0),
    .statemt_address1(grp_InversShiftRow_ByteS_fu_569_statemt_address1),
    .statemt_ce1(grp_InversShiftRow_ByteS_fu_569_statemt_ce1),
    .statemt_we1(grp_InversShiftRow_ByteS_fu_569_statemt_we1),
    .statemt_d1(grp_InversShiftRow_ByteS_fu_569_statemt_d1),
    .statemt_q1(statemt_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_AddRoundKey_InversMi_fu_548_ap_start_reg <= 1'b0;
    end else
      if((icmp_ln21_fu_594_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
        grp_AddRoundKey_InversMi_fu_548_ap_start_reg <= 1'b1;
      end else if(grp_AddRoundKey_InversMi_fu_548_ap_ready == 1'b1) begin
        grp_AddRoundKey_InversMi_fu_548_ap_start_reg <= 1'b0;
      end 
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_AddRoundKey_fu_558_ap_start_reg <= 1'b0;
    end else
      if((icmp_ln11_fu_577_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state7) & (icmp_ln21_fu_594_p2 == 1'd1)) begin
        grp_AddRoundKey_fu_558_ap_start_reg <= 1'b1;
      end else if(grp_AddRoundKey_fu_558_ap_ready == 1'b1) begin
        grp_AddRoundKey_fu_558_ap_start_reg <= 1'b0;
      end 
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_InversShiftRow_ByteS_fu_569_ap_start_reg <= 1'b0;
    end else
      if((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state5)) begin
        grp_InversShiftRow_ByteS_fu_569_ap_start_reg <= 1'b1;
      end else if(grp_InversShiftRow_ByteS_fu_569_ap_ready == 1'b1) begin
        grp_InversShiftRow_ByteS_fu_569_ap_start_reg <= 1'b0;
      end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      i_0_reg_525 <= i_reg_609;
    end else if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      i_0_reg_525 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
      if((1'b1 == ap_CS_fsm_state10) & (grp_InversShiftRow_ByteS_fu_569_ap_done == 1'b1)) begin
        i_1_reg_536 <= i_2_reg_627;
      end else if((1'b1 == ap_CS_fsm_state6) & (grp_InversShiftRow_ByteS_fu_569_ap_done == 1'b1)) begin
        i_1_reg_536 <= 4'd9;
      end  
  end


  always @(posedge ap_clk) begin
    if((icmp_ln21_fu_594_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      i_2_reg_627 <= i_2_fu_600_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state2) begin
      i_reg_609 <= i_fu_583_p2;
    end 
  end

  assign zext_ln12_fu_589_p1_temp_0 = zext_ln12_fu_589_p1 & 6'd63;
  assign zext_ln12_reg_614_temp_1 = zext_ln12_reg_614 & 6'd18446744073709551552;
  assign zext_ln12_fu_589_p1_temp_0_temp_2 = zext_ln12_fu_589_p1_temp_0 | zext_ln12_reg_614_temp_1;

  always @(posedge ap_clk) begin
    if((icmp_ln11_fu_577_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      zext_ln12_reg_614 <= zext_ln12_fu_589_p1_temp_0_temp_2;
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      grp_AddRoundKey_fu_558_n = 5'd0;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      grp_AddRoundKey_fu_558_n = 5'd10;
    end else begin
      grp_AddRoundKey_fu_558_n = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      statemt1_address0 = 64'd31;
    end else if(1'b1 == ap_CS_fsm_state27) begin
      statemt1_address0 = 64'd29;
    end else if(1'b1 == ap_CS_fsm_state26) begin
      statemt1_address0 = 64'd27;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      statemt1_address0 = 64'd25;
    end else if(1'b1 == ap_CS_fsm_state24) begin
      statemt1_address0 = 64'd23;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      statemt1_address0 = 64'd21;
    end else if(1'b1 == ap_CS_fsm_state22) begin
      statemt1_address0 = 64'd19;
    end else if(1'b1 == ap_CS_fsm_state21) begin
      statemt1_address0 = 64'd17;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt1_address0 = 64'd15;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      statemt1_address0 = 64'd13;
    end else if(1'b1 == ap_CS_fsm_state18) begin
      statemt1_address0 = 64'd11;
    end else if(1'b1 == ap_CS_fsm_state17) begin
      statemt1_address0 = 64'd9;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt1_address0 = 64'd7;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt1_address0 = 64'd5;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt1_address0 = 64'd3;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt1_address0 = 64'd0;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt1_address0 = zext_ln12_fu_589_p1;
    end else begin
      statemt1_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state28) begin
      statemt1_address1 = 64'd30;
    end else if(1'b1 == ap_CS_fsm_state27) begin
      statemt1_address1 = 64'd28;
    end else if(1'b1 == ap_CS_fsm_state26) begin
      statemt1_address1 = 64'd26;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      statemt1_address1 = 64'd24;
    end else if(1'b1 == ap_CS_fsm_state24) begin
      statemt1_address1 = 64'd22;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      statemt1_address1 = 64'd20;
    end else if(1'b1 == ap_CS_fsm_state22) begin
      statemt1_address1 = 64'd18;
    end else if(1'b1 == ap_CS_fsm_state21) begin
      statemt1_address1 = 64'd16;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt1_address1 = 64'd14;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      statemt1_address1 = 64'd12;
    end else if(1'b1 == ap_CS_fsm_state18) begin
      statemt1_address1 = 64'd10;
    end else if(1'b1 == ap_CS_fsm_state17) begin
      statemt1_address1 = 64'd8;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt1_address1 = 64'd6;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt1_address1 = 64'd4;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt1_address1 = 64'd2;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt1_address1 = 64'd1;
    end else begin
      statemt1_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt1_ce0 = 1'b1;
    end else begin
      statemt1_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt1_ce1 = 1'b1;
    end else begin
      statemt1_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt1_we0 = 1'b1;
    end else begin
      statemt1_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt1_we1 = 1'b1;
    end else begin
      statemt1_we1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      statemt_address0 = 5'd31;
    end else if(1'b1 == ap_CS_fsm_state26) begin
      statemt_address0 = 5'd29;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      statemt_address0 = 5'd27;
    end else if(1'b1 == ap_CS_fsm_state24) begin
      statemt_address0 = 5'd25;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      statemt_address0 = 5'd23;
    end else if(1'b1 == ap_CS_fsm_state22) begin
      statemt_address0 = 5'd21;
    end else if(1'b1 == ap_CS_fsm_state21) begin
      statemt_address0 = 5'd19;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_address0 = 5'd17;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      statemt_address0 = 5'd15;
    end else if(1'b1 == ap_CS_fsm_state18) begin
      statemt_address0 = 5'd13;
    end else if(1'b1 == ap_CS_fsm_state17) begin
      statemt_address0 = 5'd11;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt_address0 = 5'd9;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_address0 = 5'd7;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address0 = 5'd5;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address0 = 5'd3;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address0 = 5'd0;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = zext_ln12_reg_614;
    end else if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_address0 = grp_InversShiftRow_ByteS_fu_569_statemt_address0;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_address0 = grp_AddRoundKey_fu_558_statemt_address0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = grp_AddRoundKey_InversMi_fu_548_statemt_address0;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      statemt_address1 = 5'd30;
    end else if(1'b1 == ap_CS_fsm_state26) begin
      statemt_address1 = 5'd28;
    end else if(1'b1 == ap_CS_fsm_state25) begin
      statemt_address1 = 5'd26;
    end else if(1'b1 == ap_CS_fsm_state24) begin
      statemt_address1 = 5'd24;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      statemt_address1 = 5'd22;
    end else if(1'b1 == ap_CS_fsm_state22) begin
      statemt_address1 = 5'd20;
    end else if(1'b1 == ap_CS_fsm_state21) begin
      statemt_address1 = 5'd18;
    end else if(1'b1 == ap_CS_fsm_state20) begin
      statemt_address1 = 5'd16;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      statemt_address1 = 5'd14;
    end else if(1'b1 == ap_CS_fsm_state18) begin
      statemt_address1 = 5'd12;
    end else if(1'b1 == ap_CS_fsm_state17) begin
      statemt_address1 = 5'd10;
    end else if(1'b1 == ap_CS_fsm_state16) begin
      statemt_address1 = 5'd8;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_address1 = 5'd6;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address1 = 5'd4;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address1 = 5'd2;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address1 = 5'd1;
    end else if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_address1 = grp_InversShiftRow_ByteS_fu_569_statemt_address1;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_address1 = grp_AddRoundKey_fu_558_statemt_address1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = grp_AddRoundKey_InversMi_fu_548_statemt_address1;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state3)) begin
      statemt_ce0 = 1'b1;
    end else if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_ce0 = grp_InversShiftRow_ByteS_fu_569_statemt_ce0;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_ce0 = grp_AddRoundKey_fu_558_statemt_ce0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_ce0 = grp_AddRoundKey_InversMi_fu_548_statemt_ce0;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state26) | (1'b1 == ap_CS_fsm_state25) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state22) | (1'b1 == ap_CS_fsm_state21) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state18) | (1'b1 == ap_CS_fsm_state17) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state13)) begin
      statemt_ce1 = 1'b1;
    end else if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_ce1 = grp_InversShiftRow_ByteS_fu_569_statemt_ce1;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_ce1 = grp_AddRoundKey_fu_558_statemt_ce1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_ce1 = grp_AddRoundKey_InversMi_fu_548_statemt_ce1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_d0 = statemt1_q0;
    end else if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_d0 = grp_InversShiftRow_ByteS_fu_569_statemt_d0;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_d0 = grp_AddRoundKey_fu_558_statemt_d0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_d0 = grp_AddRoundKey_InversMi_fu_548_statemt_d0;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_d1 = grp_InversShiftRow_ByteS_fu_569_statemt_d1;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_d1 = grp_AddRoundKey_fu_558_statemt_d1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_d1 = grp_AddRoundKey_InversMi_fu_548_statemt_d1;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      statemt_we0 = 1'b1;
    end else if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_we0 = grp_InversShiftRow_ByteS_fu_569_statemt_we0;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_we0 = grp_AddRoundKey_fu_558_statemt_we0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_we0 = grp_AddRoundKey_InversMi_fu_548_statemt_we0;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state6)) begin
      statemt_we1 = grp_InversShiftRow_ByteS_fu_569_statemt_we1;
    end else if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      statemt_we1 = grp_AddRoundKey_fu_558_statemt_we1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_we1 = grp_AddRoundKey_InversMi_fu_548_statemt_we1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      word_address0 = grp_AddRoundKey_fu_558_word_address0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      word_address0 = grp_AddRoundKey_InversMi_fu_548_word_address0;
    end else begin
      word_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      word_address1 = grp_AddRoundKey_fu_558_word_address1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      word_address1 = grp_AddRoundKey_InversMi_fu_548_word_address1;
    end else begin
      word_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      word_ce0 = grp_AddRoundKey_fu_558_word_ce0;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      word_ce0 = grp_AddRoundKey_InversMi_fu_548_word_ce0;
    end else begin
      word_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state4)) begin
      word_ce1 = grp_AddRoundKey_fu_558_word_ce1;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      word_ce1 = grp_AddRoundKey_InversMi_fu_548_word_ce1;
    end else begin
      word_ce1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((icmp_ln11_fu_577_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state2;
      end
      ap_ST_fsm_state4: begin
        if((1'b1 == ap_CS_fsm_state4) & (grp_AddRoundKey_fu_558_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state5;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state6;
      end
      ap_ST_fsm_state6: begin
        if((1'b1 == ap_CS_fsm_state6) & (grp_InversShiftRow_ByteS_fu_569_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state7: begin
        if((1'b1 == ap_CS_fsm_state7) & (icmp_ln21_fu_594_p2 == 1'd1)) begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        if((1'b1 == ap_CS_fsm_state8) & (grp_AddRoundKey_InversMi_fu_548_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state9;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        if((1'b1 == ap_CS_fsm_state10) & (grp_InversShiftRow_ByteS_fu_569_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end
      end
      ap_ST_fsm_state11: begin
        if((1'b1 == ap_CS_fsm_state11) & (grp_AddRoundKey_fu_558_ap_done == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end
      end
      ap_ST_fsm_state12: begin
        ap_NS_fsm = ap_ST_fsm_state13;
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        ap_NS_fsm = ap_ST_fsm_state18;
      end
      ap_ST_fsm_state18: begin
        ap_NS_fsm = ap_ST_fsm_state19;
      end
      ap_ST_fsm_state19: begin
        ap_NS_fsm = ap_ST_fsm_state20;
      end
      ap_ST_fsm_state20: begin
        ap_NS_fsm = ap_ST_fsm_state21;
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state22;
      end
      ap_ST_fsm_state22: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state23: begin
        ap_NS_fsm = ap_ST_fsm_state24;
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state25;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state26;
      end
      ap_ST_fsm_state26: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      ap_ST_fsm_state27: begin
        ap_NS_fsm = ap_ST_fsm_state28;
      end
      ap_ST_fsm_state28: begin
        ap_NS_fsm = ap_ST_fsm_state1;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];
  assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];
  assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];
  assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];
  assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];
  assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign grp_AddRoundKey_InversMi_fu_548_ap_start = grp_AddRoundKey_InversMi_fu_548_ap_start_reg;
  assign grp_AddRoundKey_fu_558_ap_start = grp_AddRoundKey_fu_558_ap_start_reg;
  assign grp_InversShiftRow_ByteS_fu_569_ap_start = grp_InversShiftRow_ByteS_fu_569_ap_start_reg;
  assign i_2_fu_600_p2 = $signed(i_1_reg_536) + $signed(4'd15);
  assign i_fu_583_p2 = i_0_reg_525 + 6'd1;
  assign icmp_ln11_fu_577_p2 = (i_0_reg_525 == 6'd32)? 1'b1 : 1'b0;
  assign icmp_ln21_fu_594_p2 = (i_1_reg_536 == 4'd0)? 1'b1 : 1'b0;
  assign statemt1_d0 = statemt_q0;
  assign statemt1_d1 = statemt_q1;
  assign zext_ln12_fu_589_p1 = i_0_reg_525;

  always @(posedge ap_clk) begin
    zext_ln12_reg_614 <= zext_ln12_reg_614 & 63'd63;
  end


endmodule

