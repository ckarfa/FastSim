
module ByteSub_ShiftRow
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  statemt_address0,
  statemt_ce0,
  statemt_we0,
  statemt_d0,
  statemt_q0,
  statemt_address1,
  statemt_ce1,
  statemt_we1,
  statemt_d1,
  statemt_q1
);

  parameter ap_ST_fsm_state1 = 16'd1;
  parameter ap_ST_fsm_state2 = 16'd2;
  parameter ap_ST_fsm_state3 = 16'd4;
  parameter ap_ST_fsm_state4 = 16'd8;
  parameter ap_ST_fsm_state5 = 16'd16;
  parameter ap_ST_fsm_state6 = 16'd32;
  parameter ap_ST_fsm_state7 = 16'd64;
  parameter ap_ST_fsm_state8 = 16'd128;
  parameter ap_ST_fsm_state9 = 16'd256;
  parameter ap_ST_fsm_state10 = 16'd512;
  parameter ap_ST_fsm_state11 = 16'd1024;
  parameter ap_ST_fsm_state12 = 16'd2048;
  parameter ap_ST_fsm_state13 = 16'd4096;
  parameter ap_ST_fsm_state14 = 16'd8192;
  parameter ap_ST_fsm_state15 = 16'd16384;
  parameter ap_ST_fsm_state16 = 16'd32768;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  output [4:0] statemt_address0;
  output statemt_ce0;
  output statemt_we0;
  output [31:0] statemt_d0;
  input [31:0] statemt_q0;
  output [4:0] statemt_address1;
  output statemt_ce1;
  output statemt_we1;
  output [31:0] statemt_d1;
  input [31:0] statemt_q1;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [4:0] statemt_address0;
  reg statemt_ce0;
  reg statemt_we0;
  reg [31:0] statemt_d0;
  reg [4:0] statemt_address1;
  reg statemt_ce1;
  reg statemt_we1;
  reg [31:0] statemt_d1;
  reg [15:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [7:0] Sbox_address0;
  reg Sbox_ce0;
  wire [7:0] Sbox_q0;
  reg [7:0] Sbox_address1;
  reg Sbox_ce1;
  wire [7:0] Sbox_q1;
  reg [7:0] reg_338;
  wire ap_CS_fsm_state3;
  wire ap_CS_fsm_state10;
  reg [7:0] reg_342;
  wire ap_CS_fsm_state9;
  reg [7:0] reg_347;
  wire ap_CS_fsm_state4;
  reg [7:0] reg_352;
  wire [4:0] statemt_addr_21_reg_428;
  wire [4:0] statemt_addr_22_reg_433;
  wire ap_CS_fsm_state2;
  wire [4:0] statemt_addr_23_reg_448;
  wire [4:0] statemt_addr_24_reg_453;
  wire [7:0] Sbox_addr_2_gep_fu_104_p3;
  wire [7:0] Sbox_addr_3_gep_fu_113_p3;
  wire [4:0] statemt_addr_25_reg_468;
  wire [4:0] statemt_addr_26_reg_473;
  wire [7:0] Sbox_addr_4_gep_fu_140_p3;
  wire [7:0] Sbox_addr_5_gep_fu_149_p3;
  wire [4:0] statemt_addr_27_reg_488;
  wire [4:0] statemt_addr_28_reg_493;
  reg [7:0] temp_1_reg_498;
  wire ap_CS_fsm_state5;
  reg [7:0] Sbox_load_4_reg_503;
  wire [7:0] Sbox_addr_6_gep_fu_176_p3;
  wire [7:0] Sbox_addr_7_gep_fu_185_p3;
  wire [4:0] statemt_addr_29_reg_518;
  wire [4:0] statemt_addr_30_reg_523;
  reg [7:0] temp_2_reg_528;
  wire ap_CS_fsm_state6;
  reg [7:0] Sbox_load_6_reg_533;
  wire [7:0] Sbox_addr_8_gep_fu_212_p3;
  wire [7:0] Sbox_addr_9_gep_fu_221_p3;
  wire [4:0] statemt_addr_31_reg_548;
  wire [4:0] statemt_addr_32_reg_553;
  wire [4:0] statemt_addr_reg_558;
  wire ap_CS_fsm_state7;
  reg [7:0] temp_3_reg_563;
  reg [7:0] Sbox_load_8_reg_568;
  wire [7:0] Sbox_addr_10_gep_fu_256_p3;
  wire [7:0] Sbox_addr_11_gep_fu_265_p3;
  wire [4:0] statemt_addr_33_reg_583;
  reg [7:0] Sbox_load_9_reg_588;
  wire ap_CS_fsm_state8;
  reg [7:0] Sbox_load_10_reg_593;
  wire [7:0] Sbox_addr_12_gep_fu_284_p3;
  wire [7:0] Sbox_addr_13_gep_fu_293_p3;
  wire [4:0] statemt_addr_34_reg_608;
  wire [4:0] statemt_addr_35_reg_613;
  wire [7:0] Sbox_addr_14_gep_fu_320_p3;
  wire [7:0] Sbox_addr_15_gep_fu_329_p3;
  wire [31:0] Sbox_load_cast_fu_356_p1;
  wire [31:0] Sbox_load_1_cast_fu_361_p1;
  wire [31:0] Sbox_load_2_cast_fu_371_p1;
  wire [31:0] temp_cast_fu_366_p1;
  wire ap_CS_fsm_state11;
  wire [31:0] Sbox_load_4_cast_fu_380_p1;
  wire [31:0] temp_1_cast_fu_376_p1;
  wire ap_CS_fsm_state12;
  wire [31:0] Sbox_load_6_cast_fu_388_p1;
  wire [31:0] temp_2_cast_fu_384_p1;
  wire ap_CS_fsm_state13;
  wire [31:0] Sbox_load_8_cast_fu_392_p1;
  wire [31:0] Sbox_load_9_cast_fu_396_p1;
  wire ap_CS_fsm_state14;
  wire [31:0] Sbox_load_10_cast_fu_404_p1;
  wire [31:0] temp_3_cast_fu_400_p1;
  wire ap_CS_fsm_state15;
  wire [31:0] Sbox_load_11_cast_fu_408_p1;
  wire [31:0] Sbox_load_12_cast_fu_413_p1;
  wire ap_CS_fsm_state16;
  wire [31:0] Sbox_load_13_cast_fu_418_p1;
  wire [31:0] Sbox_load_14_cast_fu_423_p1;
  reg [15:0] ap_NS_fsm;

  initial begin
    #0 ap_CS_fsm = 16'd1;
  end


  KeySchedule_Sbox
  #(
    .DataWidth(8),
    .AddressRange(256),
    .AddressWidth(8)
  )
  Sbox_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(Sbox_address0),
    .ce0(Sbox_ce0),
    .q0(Sbox_q0),
    .address1(Sbox_address1),
    .ce1(Sbox_ce1),
    .q1(Sbox_q1)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      reg_342 <= Sbox_q0;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      reg_342 <= Sbox_q1;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      reg_347 <= Sbox_q1;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      reg_347 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state8) begin
      Sbox_load_10_reg_593 <= Sbox_q1;
      Sbox_load_9_reg_588 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      Sbox_load_4_reg_503 <= Sbox_q1;
      temp_1_reg_498 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state6) begin
      Sbox_load_6_reg_533 <= Sbox_q1;
      temp_2_reg_528 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_load_8_reg_568 <= Sbox_q1;
      temp_3_reg_563 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state10)) begin
      reg_338 <= Sbox_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state4)) begin
      reg_352 <= Sbox_q1;
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      Sbox_address0 = Sbox_addr_14_gep_fu_320_p3;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      Sbox_address0 = Sbox_addr_12_gep_fu_284_p3;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_address0 = Sbox_addr_10_gep_fu_256_p3;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      Sbox_address0 = Sbox_addr_8_gep_fu_212_p3;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      Sbox_address0 = Sbox_addr_6_gep_fu_176_p3;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      Sbox_address0 = Sbox_addr_4_gep_fu_140_p3;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      Sbox_address0 = Sbox_addr_2_gep_fu_104_p3;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      Sbox_address0 = statemt_q0;
    end else begin
      Sbox_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      Sbox_address1 = Sbox_addr_15_gep_fu_329_p3;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      Sbox_address1 = Sbox_addr_13_gep_fu_293_p3;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      Sbox_address1 = Sbox_addr_11_gep_fu_265_p3;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      Sbox_address1 = Sbox_addr_9_gep_fu_221_p3;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      Sbox_address1 = Sbox_addr_7_gep_fu_185_p3;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      Sbox_address1 = Sbox_addr_5_gep_fu_149_p3;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      Sbox_address1 = Sbox_addr_3_gep_fu_113_p3;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      Sbox_address1 = statemt_q1;
    end else begin
      Sbox_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state8)) begin
      Sbox_ce0 = 1'b1;
    end else begin
      Sbox_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state8)) begin
      Sbox_ce1 = 1'b1;
    end else begin
      Sbox_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_start) & (1'b1 == ap_CS_fsm_state1) | (1'b1 == ap_CS_fsm_state16)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((1'b0 == ap_start) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_address0 = statemt_addr_34_reg_608;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_address0 = statemt_addr_reg_558;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address0 = statemt_addr_31_reg_548;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address0 = statemt_addr_29_reg_518;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address0 = statemt_addr_27_reg_488;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_address0 = statemt_addr_25_reg_468;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_address0 = statemt_addr_23_reg_448;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_address0 = statemt_addr_21_reg_428;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address0 = 32'd8;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address0 = 32'd0;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      statemt_address0 = 32'd11;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address0 = 32'd3;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address0 = 32'd6;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address0 = 32'd2;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address0 = 32'd9;
    end else if(1'b1 == ap_CS_fsm_state1) begin
      statemt_address0 = 32'd1;
    end else begin
      statemt_address0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_address1 = statemt_addr_35_reg_613;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_address1 = statemt_addr_33_reg_583;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_address1 = statemt_addr_32_reg_553;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_address1 = statemt_addr_30_reg_523;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_address1 = statemt_addr_28_reg_493;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_address1 = statemt_addr_26_reg_473;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_address1 = statemt_addr_24_reg_453;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_address1 = statemt_addr_22_reg_433;
    end else if(1'b1 == ap_CS_fsm_state8) begin
      statemt_address1 = 32'd12;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      statemt_address1 = 32'd4;
    end else if(1'b1 == ap_CS_fsm_state6) begin
      statemt_address1 = 32'd7;
    end else if(1'b1 == ap_CS_fsm_state5) begin
      statemt_address1 = 32'd15;
    end else if(1'b1 == ap_CS_fsm_state4) begin
      statemt_address1 = 32'd14;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      statemt_address1 = 32'd10;
    end else if(1'b1 == ap_CS_fsm_state2) begin
      statemt_address1 = 32'd13;
    end else if(1'b1 == ap_CS_fsm_state1) begin
      statemt_address1 = 32'd5;
    end else begin
      statemt_address1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state16)) begin
      statemt_ce0 = 1'b1;
    end else begin
      statemt_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state3) | (1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state4) | (1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1) | (1'b1 == ap_CS_fsm_state2) | (1'b1 == ap_CS_fsm_state5) | (1'b1 == ap_CS_fsm_state6) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state16)) begin
      statemt_ce1 = 1'b1;
    end else begin
      statemt_ce1 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_d0 = Sbox_load_13_cast_fu_418_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_d0 = Sbox_load_11_cast_fu_408_p1;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d0 = Sbox_load_10_cast_fu_404_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d0 = Sbox_load_8_cast_fu_392_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_d0 = Sbox_load_6_cast_fu_388_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_d0 = Sbox_load_4_cast_fu_380_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_d0 = Sbox_load_2_cast_fu_371_p1;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_d0 = Sbox_load_cast_fu_356_p1;
    end else begin
      statemt_d0 = 'bx;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state16) begin
      statemt_d1 = Sbox_load_14_cast_fu_423_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      statemt_d1 = Sbox_load_12_cast_fu_413_p1;
    end else if(1'b1 == ap_CS_fsm_state14) begin
      statemt_d1 = temp_3_cast_fu_400_p1;
    end else if(1'b1 == ap_CS_fsm_state13) begin
      statemt_d1 = Sbox_load_9_cast_fu_396_p1;
    end else if(1'b1 == ap_CS_fsm_state12) begin
      statemt_d1 = temp_2_cast_fu_384_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      statemt_d1 = temp_1_cast_fu_376_p1;
    end else if(1'b1 == ap_CS_fsm_state10) begin
      statemt_d1 = temp_cast_fu_366_p1;
    end else if(1'b1 == ap_CS_fsm_state9) begin
      statemt_d1 = Sbox_load_1_cast_fu_361_p1;
    end else begin
      statemt_d1 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state16)) begin
      statemt_we0 = 1'b1;
    end else begin
      statemt_we0 = 1'b0;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state10) | (1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state14) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state16)) begin
      statemt_we1 = 1'b1;
    end else begin
      statemt_we1 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        ap_NS_fsm = ap_ST_fsm_state3;
      end
      ap_ST_fsm_state3: begin
        ap_NS_fsm = ap_ST_fsm_state4;
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state6;
      end
      ap_ST_fsm_state6: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state7: begin
        ap_NS_fsm = ap_ST_fsm_state8;
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state10;
      end
      ap_ST_fsm_state10: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state11: begin
        ap_NS_fsm = ap_ST_fsm_state12;
      end
      ap_ST_fsm_state12: begin
        ap_NS_fsm = ap_ST_fsm_state13;
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state14;
      end
      ap_ST_fsm_state14: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state15: begin
        ap_NS_fsm = ap_ST_fsm_state16;
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state1;
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign Sbox_addr_10_gep_fu_256_p3 = statemt_q0;
  assign Sbox_addr_11_gep_fu_265_p3 = statemt_q1;
  assign Sbox_addr_12_gep_fu_284_p3 = statemt_q0;
  assign Sbox_addr_13_gep_fu_293_p3 = statemt_q1;
  assign Sbox_addr_14_gep_fu_320_p3 = statemt_q0;
  assign Sbox_addr_15_gep_fu_329_p3 = statemt_q1;
  assign Sbox_addr_2_gep_fu_104_p3 = statemt_q0;
  assign Sbox_addr_3_gep_fu_113_p3 = statemt_q1;
  assign Sbox_addr_4_gep_fu_140_p3 = statemt_q0;
  assign Sbox_addr_5_gep_fu_149_p3 = statemt_q1;
  assign Sbox_addr_6_gep_fu_176_p3 = statemt_q0;
  assign Sbox_addr_7_gep_fu_185_p3 = statemt_q1;
  assign Sbox_addr_8_gep_fu_212_p3 = statemt_q0;
  assign Sbox_addr_9_gep_fu_221_p3 = statemt_q1;
  assign Sbox_load_10_cast_fu_404_p1 = Sbox_load_10_reg_593;
  assign Sbox_load_11_cast_fu_408_p1 = reg_342;
  assign Sbox_load_12_cast_fu_413_p1 = reg_347;
  assign Sbox_load_13_cast_fu_418_p1 = reg_338;
  assign Sbox_load_14_cast_fu_423_p1 = reg_352;
  assign Sbox_load_1_cast_fu_361_p1 = reg_347;
  assign Sbox_load_2_cast_fu_371_p1 = reg_352;
  assign Sbox_load_4_cast_fu_380_p1 = Sbox_load_4_reg_503;
  assign Sbox_load_6_cast_fu_388_p1 = Sbox_load_6_reg_533;
  assign Sbox_load_8_cast_fu_392_p1 = Sbox_load_8_reg_568;
  assign Sbox_load_9_cast_fu_396_p1 = Sbox_load_9_reg_588;
  assign Sbox_load_cast_fu_356_p1 = reg_342;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign statemt_addr_21_reg_428 = 32'd1;
  assign statemt_addr_22_reg_433 = 32'd5;
  assign statemt_addr_23_reg_448 = 32'd9;
  assign statemt_addr_24_reg_453 = 32'd13;
  assign statemt_addr_25_reg_468 = 32'd2;
  assign statemt_addr_26_reg_473 = 32'd10;
  assign statemt_addr_27_reg_488 = 32'd6;
  assign statemt_addr_28_reg_493 = 32'd14;
  assign statemt_addr_29_reg_518 = 32'd3;
  assign statemt_addr_30_reg_523 = 32'd15;
  assign statemt_addr_31_reg_548 = 32'd11;
  assign statemt_addr_32_reg_553 = 32'd7;
  assign statemt_addr_33_reg_583 = 32'd4;
  assign statemt_addr_34_reg_608 = 32'd8;
  assign statemt_addr_35_reg_613 = 32'd12;
  assign statemt_addr_reg_558 = 32'd0;
  assign temp_1_cast_fu_376_p1 = temp_1_reg_498;
  assign temp_2_cast_fu_384_p1 = temp_2_reg_528;
  assign temp_3_cast_fu_400_p1 = temp_3_reg_563;
  assign temp_cast_fu_366_p1 = reg_338;

endmodule

