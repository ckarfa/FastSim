
module insertion_cell_sort
(
  in_V_dout,
  in_V_empty_n,
  in_V_read,
  out_V_din,
  out_V_full_n,
  out_V_write,
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_ready,
  ap_idle
);

  input [31:0] in_V_dout;
  input in_V_empty_n;
  output in_V_read;
  output [31:0] out_V_din;
  input out_V_full_n;
  output out_V_write;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_ready;
  output ap_idle;
  wire cell0_U0_ap_start;
  wire cell0_U0_ap_done;
  wire cell0_U0_ap_continue;
  wire cell0_U0_ap_idle;
  wire cell0_U0_ap_ready;
  wire cell0_U0_start_out;
  wire cell0_U0_start_write;
  wire cell0_U0_in_V_read;
  wire [31:0] cell0_U0_out_V_din;
  wire cell0_U0_out_V_write;
  wire cell1_U0_ap_start;
  wire cell1_U0_ap_done;
  wire cell1_U0_ap_continue;
  wire cell1_U0_ap_idle;
  wire cell1_U0_ap_ready;
  wire cell1_U0_start_out;
  wire cell1_U0_start_write;
  wire cell1_U0_in_V_read;
  wire [31:0] cell1_U0_out_V_din;
  wire cell1_U0_out_V_write;
  wire cell2_U0_ap_start;
  wire cell2_U0_ap_done;
  wire cell2_U0_ap_continue;
  wire cell2_U0_ap_idle;
  wire cell2_U0_ap_ready;
  wire cell2_U0_start_out;
  wire cell2_U0_start_write;
  wire cell2_U0_in_V_read;
  wire [31:0] cell2_U0_out_V_din;
  wire cell2_U0_out_V_write;
  wire cell3_U0_ap_start;
  wire cell3_U0_ap_done;
  wire cell3_U0_ap_continue;
  wire cell3_U0_ap_idle;
  wire cell3_U0_ap_ready;
  wire cell3_U0_start_out;
  wire cell3_U0_start_write;
  wire cell3_U0_in_V_read;
  wire [31:0] cell3_U0_out_V_din;
  wire cell3_U0_out_V_write;
  wire cell4_U0_ap_start;
  wire cell4_U0_ap_done;
  wire cell4_U0_ap_continue;
  wire cell4_U0_ap_idle;
  wire cell4_U0_ap_ready;
  wire cell4_U0_start_out;
  wire cell4_U0_start_write;
  wire cell4_U0_in_V_read;
  wire [31:0] cell4_U0_out_V_din;
  wire cell4_U0_out_V_write;
  wire cell5_U0_ap_start;
  wire cell5_U0_ap_done;
  wire cell5_U0_ap_continue;
  wire cell5_U0_ap_idle;
  wire cell5_U0_ap_ready;
  wire cell5_U0_start_out;
  wire cell5_U0_start_write;
  wire cell5_U0_in_V_read;
  wire [31:0] cell5_U0_out_V_din;
  wire cell5_U0_out_V_write;
  wire cell6_U0_ap_start;
  wire cell6_U0_ap_done;
  wire cell6_U0_ap_continue;
  wire cell6_U0_ap_idle;
  wire cell6_U0_ap_ready;
  wire cell6_U0_start_out;
  wire cell6_U0_start_write;
  wire cell6_U0_in_V_read;
  wire [31:0] cell6_U0_out_V_din;
  wire cell6_U0_out_V_write;
  wire cell7_U0_ap_start;
  wire cell7_U0_ap_done;
  wire cell7_U0_ap_continue;
  wire cell7_U0_ap_idle;
  wire cell7_U0_ap_ready;
  wire cell7_U0_in_V_read;
  wire [31:0] cell7_U0_out_V_din;
  wire cell7_U0_out_V_write;
  wire ap_sync_continue;
  wire out1_V_full_n;
  wire [31:0] out1_V_dout;
  wire out1_V_empty_n;
  wire out2_V_full_n;
  wire [31:0] out2_V_dout;
  wire out2_V_empty_n;
  wire out3_V_full_n;
  wire [31:0] out3_V_dout;
  wire out3_V_empty_n;
  wire out4_V_full_n;
  wire [31:0] out4_V_dout;
  wire out4_V_empty_n;
  wire out5_V_full_n;
  wire [31:0] out5_V_dout;
  wire out5_V_empty_n;
  wire out6_V_full_n;
  wire [31:0] out6_V_dout;
  wire out6_V_empty_n;
  wire out7_V_full_n;
  wire [31:0] out7_V_dout;
  wire out7_V_empty_n;
  wire ap_sync_done;
  wire ap_sync_ready;
  wire [0:0] start_for_cell1_U0_din;
  wire start_for_cell1_U0_full_n;
  wire [0:0] start_for_cell1_U0_dout;
  wire start_for_cell1_U0_empty_n;
  wire [0:0] start_for_cell2_U0_din;
  wire start_for_cell2_U0_full_n;
  wire [0:0] start_for_cell2_U0_dout;
  wire start_for_cell2_U0_empty_n;
  wire [0:0] start_for_cell3_U0_din;
  wire start_for_cell3_U0_full_n;
  wire [0:0] start_for_cell3_U0_dout;
  wire start_for_cell3_U0_empty_n;
  wire [0:0] start_for_cell4_U0_din;
  wire start_for_cell4_U0_full_n;
  wire [0:0] start_for_cell4_U0_dout;
  wire start_for_cell4_U0_empty_n;
  wire [0:0] start_for_cell5_U0_din;
  wire start_for_cell5_U0_full_n;
  wire [0:0] start_for_cell5_U0_dout;
  wire start_for_cell5_U0_empty_n;
  wire [0:0] start_for_cell6_U0_din;
  wire start_for_cell6_U0_full_n;
  wire [0:0] start_for_cell6_U0_dout;
  wire start_for_cell6_U0_empty_n;
  wire [0:0] start_for_cell7_U0_din;
  wire start_for_cell7_U0_full_n;
  wire [0:0] start_for_cell7_U0_dout;
  wire start_for_cell7_U0_empty_n;
  wire cell7_U0_start_full_n;
  wire cell7_U0_start_write;

  cell0
  cell0_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell0_U0_ap_start),
    .start_full_n(start_for_cell1_U0_full_n),
    .ap_done(cell0_U0_ap_done),
    .ap_continue(cell0_U0_ap_continue),
    .ap_idle(cell0_U0_ap_idle),
    .ap_ready(cell0_U0_ap_ready),
    .start_out(cell0_U0_start_out),
    .start_write(cell0_U0_start_write),
    .in_V_dout(in_V_dout),
    .in_V_empty_n(in_V_empty_n),
    .in_V_read(cell0_U0_in_V_read),
    .out_V_din(cell0_U0_out_V_din),
    .out_V_full_n(out1_V_full_n),
    .out_V_write(cell0_U0_out_V_write)
  );


  cell1
  cell1_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell1_U0_ap_start),
    .start_full_n(start_for_cell2_U0_full_n),
    .ap_done(cell1_U0_ap_done),
    .ap_continue(cell1_U0_ap_continue),
    .ap_idle(cell1_U0_ap_idle),
    .ap_ready(cell1_U0_ap_ready),
    .start_out(cell1_U0_start_out),
    .start_write(cell1_U0_start_write),
    .in_V_dout(out1_V_dout),
    .in_V_empty_n(out1_V_empty_n),
    .in_V_read(cell1_U0_in_V_read),
    .out_V_din(cell1_U0_out_V_din),
    .out_V_full_n(out2_V_full_n),
    .out_V_write(cell1_U0_out_V_write)
  );


  cell2
  cell2_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell2_U0_ap_start),
    .start_full_n(start_for_cell3_U0_full_n),
    .ap_done(cell2_U0_ap_done),
    .ap_continue(cell2_U0_ap_continue),
    .ap_idle(cell2_U0_ap_idle),
    .ap_ready(cell2_U0_ap_ready),
    .start_out(cell2_U0_start_out),
    .start_write(cell2_U0_start_write),
    .in_V_dout(out2_V_dout),
    .in_V_empty_n(out2_V_empty_n),
    .in_V_read(cell2_U0_in_V_read),
    .out_V_din(cell2_U0_out_V_din),
    .out_V_full_n(out3_V_full_n),
    .out_V_write(cell2_U0_out_V_write)
  );


  cell3
  cell3_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell3_U0_ap_start),
    .start_full_n(start_for_cell4_U0_full_n),
    .ap_done(cell3_U0_ap_done),
    .ap_continue(cell3_U0_ap_continue),
    .ap_idle(cell3_U0_ap_idle),
    .ap_ready(cell3_U0_ap_ready),
    .start_out(cell3_U0_start_out),
    .start_write(cell3_U0_start_write),
    .in_V_dout(out3_V_dout),
    .in_V_empty_n(out3_V_empty_n),
    .in_V_read(cell3_U0_in_V_read),
    .out_V_din(cell3_U0_out_V_din),
    .out_V_full_n(out4_V_full_n),
    .out_V_write(cell3_U0_out_V_write)
  );


  cell4
  cell4_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell4_U0_ap_start),
    .start_full_n(start_for_cell5_U0_full_n),
    .ap_done(cell4_U0_ap_done),
    .ap_continue(cell4_U0_ap_continue),
    .ap_idle(cell4_U0_ap_idle),
    .ap_ready(cell4_U0_ap_ready),
    .start_out(cell4_U0_start_out),
    .start_write(cell4_U0_start_write),
    .in_V_dout(out4_V_dout),
    .in_V_empty_n(out4_V_empty_n),
    .in_V_read(cell4_U0_in_V_read),
    .out_V_din(cell4_U0_out_V_din),
    .out_V_full_n(out5_V_full_n),
    .out_V_write(cell4_U0_out_V_write)
  );


  cell5
  cell5_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell5_U0_ap_start),
    .start_full_n(start_for_cell6_U0_full_n),
    .ap_done(cell5_U0_ap_done),
    .ap_continue(cell5_U0_ap_continue),
    .ap_idle(cell5_U0_ap_idle),
    .ap_ready(cell5_U0_ap_ready),
    .start_out(cell5_U0_start_out),
    .start_write(cell5_U0_start_write),
    .in_V_dout(out5_V_dout),
    .in_V_empty_n(out5_V_empty_n),
    .in_V_read(cell5_U0_in_V_read),
    .out_V_din(cell5_U0_out_V_din),
    .out_V_full_n(out6_V_full_n),
    .out_V_write(cell5_U0_out_V_write)
  );


  cell6
  cell6_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell6_U0_ap_start),
    .start_full_n(start_for_cell7_U0_full_n),
    .ap_done(cell6_U0_ap_done),
    .ap_continue(cell6_U0_ap_continue),
    .ap_idle(cell6_U0_ap_idle),
    .ap_ready(cell6_U0_ap_ready),
    .start_out(cell6_U0_start_out),
    .start_write(cell6_U0_start_write),
    .in_V_dout(out6_V_dout),
    .in_V_empty_n(out6_V_empty_n),
    .in_V_read(cell6_U0_in_V_read),
    .out_V_din(cell6_U0_out_V_din),
    .out_V_full_n(out7_V_full_n),
    .out_V_write(cell6_U0_out_V_write)
  );


  cell7
  cell7_U0
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(cell7_U0_ap_start),
    .ap_done(cell7_U0_ap_done),
    .ap_continue(cell7_U0_ap_continue),
    .ap_idle(cell7_U0_ap_idle),
    .ap_ready(cell7_U0_ap_ready),
    .in_V_dout(out7_V_dout),
    .in_V_empty_n(out7_V_empty_n),
    .in_V_read(cell7_U0_in_V_read),
    .out_V_din(cell7_U0_out_V_din),
    .out_V_full_n(out_V_full_n),
    .out_V_write(cell7_U0_out_V_write)
  );


  fifo_w32_d2_A
  out1_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell0_U0_out_V_din),
    .if_full_n(out1_V_full_n),
    .if_write(cell0_U0_out_V_write),
    .if_dout(out1_V_dout),
    .if_empty_n(out1_V_empty_n),
    .if_read(cell1_U0_in_V_read)
  );


  fifo_w32_d2_A
  out2_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell1_U0_out_V_din),
    .if_full_n(out2_V_full_n),
    .if_write(cell1_U0_out_V_write),
    .if_dout(out2_V_dout),
    .if_empty_n(out2_V_empty_n),
    .if_read(cell2_U0_in_V_read)
  );


  fifo_w32_d2_A
  out3_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell2_U0_out_V_din),
    .if_full_n(out3_V_full_n),
    .if_write(cell2_U0_out_V_write),
    .if_dout(out3_V_dout),
    .if_empty_n(out3_V_empty_n),
    .if_read(cell3_U0_in_V_read)
  );


  fifo_w32_d2_A
  out4_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell3_U0_out_V_din),
    .if_full_n(out4_V_full_n),
    .if_write(cell3_U0_out_V_write),
    .if_dout(out4_V_dout),
    .if_empty_n(out4_V_empty_n),
    .if_read(cell4_U0_in_V_read)
  );


  fifo_w32_d2_A
  out5_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell4_U0_out_V_din),
    .if_full_n(out5_V_full_n),
    .if_write(cell4_U0_out_V_write),
    .if_dout(out5_V_dout),
    .if_empty_n(out5_V_empty_n),
    .if_read(cell5_U0_in_V_read)
  );


  fifo_w32_d2_A
  out6_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell5_U0_out_V_din),
    .if_full_n(out6_V_full_n),
    .if_write(cell5_U0_out_V_write),
    .if_dout(out6_V_dout),
    .if_empty_n(out6_V_empty_n),
    .if_read(cell6_U0_in_V_read)
  );


  fifo_w32_d2_A
  out7_V_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(cell6_U0_out_V_din),
    .if_full_n(out7_V_full_n),
    .if_write(cell6_U0_out_V_write),
    .if_dout(out7_V_dout),
    .if_empty_n(out7_V_empty_n),
    .if_read(cell7_U0_in_V_read)
  );


  start_for_cell1_U0
  start_for_cell1_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell1_U0_din),
    .if_full_n(start_for_cell1_U0_full_n),
    .if_write(cell0_U0_start_write),
    .if_dout(start_for_cell1_U0_dout),
    .if_empty_n(start_for_cell1_U0_empty_n),
    .if_read(cell1_U0_ap_ready)
  );


  start_for_cell2_U0
  start_for_cell2_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell2_U0_din),
    .if_full_n(start_for_cell2_U0_full_n),
    .if_write(cell1_U0_start_write),
    .if_dout(start_for_cell2_U0_dout),
    .if_empty_n(start_for_cell2_U0_empty_n),
    .if_read(cell2_U0_ap_ready)
  );


  start_for_cell3_U0
  start_for_cell3_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell3_U0_din),
    .if_full_n(start_for_cell3_U0_full_n),
    .if_write(cell2_U0_start_write),
    .if_dout(start_for_cell3_U0_dout),
    .if_empty_n(start_for_cell3_U0_empty_n),
    .if_read(cell3_U0_ap_ready)
  );


  start_for_cell4_U0
  start_for_cell4_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell4_U0_din),
    .if_full_n(start_for_cell4_U0_full_n),
    .if_write(cell3_U0_start_write),
    .if_dout(start_for_cell4_U0_dout),
    .if_empty_n(start_for_cell4_U0_empty_n),
    .if_read(cell4_U0_ap_ready)
  );


  start_for_cell5_U0
  start_for_cell5_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell5_U0_din),
    .if_full_n(start_for_cell5_U0_full_n),
    .if_write(cell4_U0_start_write),
    .if_dout(start_for_cell5_U0_dout),
    .if_empty_n(start_for_cell5_U0_empty_n),
    .if_read(cell5_U0_ap_ready)
  );


  start_for_cell6_U0
  start_for_cell6_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell6_U0_din),
    .if_full_n(start_for_cell6_U0_full_n),
    .if_write(cell5_U0_start_write),
    .if_dout(start_for_cell6_U0_dout),
    .if_empty_n(start_for_cell6_U0_empty_n),
    .if_read(cell6_U0_ap_ready)
  );


  start_for_cell7_U0
  start_for_cell7_U0_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .if_read_ce(1'b1),
    .if_write_ce(1'b1),
    .if_din(start_for_cell7_U0_din),
    .if_full_n(start_for_cell7_U0_full_n),
    .if_write(cell6_U0_start_write),
    .if_dout(start_for_cell7_U0_dout),
    .if_empty_n(start_for_cell7_U0_empty_n),
    .if_read(cell7_U0_ap_ready)
  );

  assign ap_done = cell7_U0_ap_done;
  assign ap_idle = cell7_U0_ap_idle & cell6_U0_ap_idle & cell5_U0_ap_idle & cell4_U0_ap_idle & cell3_U0_ap_idle & cell2_U0_ap_idle & cell1_U0_ap_idle & cell0_U0_ap_idle;
  assign ap_ready = cell0_U0_ap_ready;
  assign ap_sync_continue = 1'b1;
  assign ap_sync_done = cell7_U0_ap_done;
  assign ap_sync_ready = cell0_U0_ap_ready;
  assign cell0_U0_ap_continue = 1'b1;
  assign cell0_U0_ap_start = ap_start;
  assign cell1_U0_ap_continue = 1'b1;
  assign cell1_U0_ap_start = start_for_cell1_U0_empty_n;
  assign cell2_U0_ap_continue = 1'b1;
  assign cell2_U0_ap_start = start_for_cell2_U0_empty_n;
  assign cell3_U0_ap_continue = 1'b1;
  assign cell3_U0_ap_start = start_for_cell3_U0_empty_n;
  assign cell4_U0_ap_continue = 1'b1;
  assign cell4_U0_ap_start = start_for_cell4_U0_empty_n;
  assign cell5_U0_ap_continue = 1'b1;
  assign cell5_U0_ap_start = start_for_cell5_U0_empty_n;
  assign cell6_U0_ap_continue = 1'b1;
  assign cell6_U0_ap_start = start_for_cell6_U0_empty_n;
  assign cell7_U0_ap_continue = 1'b1;
  assign cell7_U0_ap_start = start_for_cell7_U0_empty_n;
  assign cell7_U0_start_full_n = 1'b1;
  assign cell7_U0_start_write = 1'b0;
  assign in_V_read = cell0_U0_in_V_read;
  assign out_V_din = cell7_U0_out_V_din;
  assign out_V_write = cell7_U0_out_V_write;
  assign start_for_cell1_U0_din = 1'b1;
  assign start_for_cell2_U0_din = 1'b1;
  assign start_for_cell3_U0_din = 1'b1;
  assign start_for_cell4_U0_din = 1'b1;
  assign start_for_cell5_U0_din = 1'b1;
  assign start_for_cell6_U0_din = 1'b1;
  assign start_for_cell7_U0_din = 1'b1;

endmodule

