
module shiftingcidi
(
  ap_clk,
  ap_rst,
  ap_start,
  ap_done,
  ap_idle,
  ap_ready,
  C,
  D,
  L,
  R,
  ap_return
);

  parameter ap_ST_fsm_state1 = 67'd1;
  parameter ap_ST_fsm_state2 = 67'd2;
  parameter ap_ST_fsm_state3 = 67'd4;
  parameter ap_ST_fsm_state4 = 67'd8;
  parameter ap_ST_fsm_state5 = 67'd16;
  parameter ap_ST_fsm_state6 = 67'd32;
  parameter ap_ST_fsm_state7 = 67'd64;
  parameter ap_ST_fsm_state8 = 67'd128;
  parameter ap_ST_fsm_state9 = 67'd256;
  parameter ap_ST_fsm_state10 = 67'd512;
  parameter ap_ST_fsm_state11 = 67'd1024;
  parameter ap_ST_fsm_state12 = 67'd2048;
  parameter ap_ST_fsm_state13 = 67'd4096;
  parameter ap_ST_fsm_state14 = 67'd8192;
  parameter ap_ST_fsm_state15 = 67'd16384;
  parameter ap_ST_fsm_state16 = 67'd32768;
  parameter ap_ST_fsm_state17 = 67'd65536;
  parameter ap_ST_fsm_state18 = 67'd131072;
  parameter ap_ST_fsm_state19 = 67'd262144;
  parameter ap_ST_fsm_state20 = 67'd524288;
  parameter ap_ST_fsm_state21 = 67'd1048576;
  parameter ap_ST_fsm_state22 = 67'd2097152;
  parameter ap_ST_fsm_state23 = 67'd4194304;
  parameter ap_ST_fsm_state24 = 67'd8388608;
  parameter ap_ST_fsm_state25 = 67'd16777216;
  parameter ap_ST_fsm_state26 = 67'd33554432;
  parameter ap_ST_fsm_state27 = 67'd67108864;
  parameter ap_ST_fsm_state28 = 67'd134217728;
  parameter ap_ST_fsm_state29 = 67'd268435456;
  parameter ap_ST_fsm_state30 = 67'd536870912;
  parameter ap_ST_fsm_state31 = 67'd1073741824;
  parameter ap_ST_fsm_state32 = 67'd2147483648;
  parameter ap_ST_fsm_state33 = 67'd4294967296;
  parameter ap_ST_fsm_state34 = 67'd8589934592;
  parameter ap_ST_fsm_state35 = 67'd17179869184;
  parameter ap_ST_fsm_state36 = 67'd34359738368;
  parameter ap_ST_fsm_state37 = 67'd68719476736;
  parameter ap_ST_fsm_state38 = 67'd137438953472;
  parameter ap_ST_fsm_state39 = 67'd274877906944;
  parameter ap_ST_fsm_state40 = 67'd549755813888;
  parameter ap_ST_fsm_state41 = 67'd1099511627776;
  parameter ap_ST_fsm_state42 = 67'd2199023255552;
  parameter ap_ST_fsm_state43 = 67'd4398046511104;
  parameter ap_ST_fsm_state44 = 67'd8796093022208;
  parameter ap_ST_fsm_state45 = 67'd17592186044416;
  parameter ap_ST_fsm_state46 = 67'd35184372088832;
  parameter ap_ST_fsm_state47 = 67'd70368744177664;
  parameter ap_ST_fsm_state48 = 67'd140737488355328;
  parameter ap_ST_fsm_state49 = 67'd281474976710656;
  parameter ap_ST_fsm_state50 = 67'd562949953421312;
  parameter ap_ST_fsm_state51 = 67'd1125899906842624;
  parameter ap_ST_fsm_state52 = 67'd2251799813685248;
  parameter ap_ST_fsm_state53 = 67'd4503599627370496;
  parameter ap_ST_fsm_state54 = 67'd9007199254740992;
  parameter ap_ST_fsm_state55 = 67'd18014398509481984;
  parameter ap_ST_fsm_state56 = 67'd36028797018963968;
  parameter ap_ST_fsm_state57 = 67'd72057594037927936;
  parameter ap_ST_fsm_state58 = 67'd144115188075855872;
  parameter ap_ST_fsm_state59 = 67'd288230376151711744;
  parameter ap_ST_fsm_state60 = 67'd576460752303423488;
  parameter ap_ST_fsm_state61 = 67'd1152921504606846976;
  parameter ap_ST_fsm_state62 = 67'd2305843009213693952;
  parameter ap_ST_fsm_state63 = 67'd4611686018427387904;
  parameter ap_ST_fsm_state64 = 67'd9223372036854775808;
  parameter ap_ST_fsm_state65 = 67'd18446744073709551616;
  parameter ap_ST_fsm_state66 = 67'd36893488147419103232;
  parameter ap_ST_fsm_state67 = 67'd73786976294838206464;
  input ap_clk;
  input ap_rst;
  input ap_start;
  output ap_done;
  output ap_idle;
  output ap_ready;
  input [27:0] C;
  input [27:0] D;
  input [31:0] L;
  input [31:0] R;
  output [63:0] ap_return;
  reg ap_done;
  reg ap_idle;
  reg ap_ready;
  reg [63:0] ap_return;
  reg [66:0] ap_CS_fsm;
  wire ap_CS_fsm_state1;
  reg [5:0] PC2_address0;
  reg PC2_ce0;
  wire [5:0] PC2_q0;
  reg [3:0] sub_key_address0;
  reg sub_key_ce0;
  reg sub_key_we0;
  reg [63:0] sub_key_d0;
  wire [63:0] sub_key_q0;
  reg [5:0] reg_1192;
  wire ap_CS_fsm_state4;
  wire ap_CS_fsm_state8;
  wire ap_CS_fsm_state12;
  wire ap_CS_fsm_state16;
  wire ap_CS_fsm_state20;
  wire ap_CS_fsm_state24;
  wire ap_CS_fsm_state28;
  wire ap_CS_fsm_state32;
  wire ap_CS_fsm_state36;
  wire ap_CS_fsm_state40;
  wire ap_CS_fsm_state44;
  wire ap_CS_fsm_state48;
  wire ap_CS_fsm_state52;
  wire ap_CS_fsm_state56;
  wire ap_CS_fsm_state60;
  wire ap_CS_fsm_state64;
  wire [27:0] or_ln_fu_1214_p3;
  wire ap_CS_fsm_state2;
  wire [0:0] ap_phi_mux_j_0_0_phi_fu_304_p4;
  wire [27:0] or_ln1_fu_1234_p3;
  wire [55:0] tmp_2_fu_1242_p3;
  reg [55:0] tmp_2_reg_2800;
  wire [5:0] add_ln121_fu_1256_p2;
  reg [5:0] add_ln121_reg_2808;
  wire ap_CS_fsm_state3;
  wire [0:0] icmp_ln121_fu_1250_p2;
  wire [62:0] trunc_ln125_1_fu_1267_p1;
  reg [62:0] trunc_ln125_1_reg_2818;
  wire [63:0] or_ln2_fu_1284_p3;
  wire ap_CS_fsm_state5;
  wire [27:0] or_ln111_1_fu_1303_p3;
  wire ap_CS_fsm_state6;
  wire [0:0] ap_phi_mux_j_0_1_phi_fu_361_p4;
  wire [27:0] or_ln113_1_fu_1323_p3;
  wire [55:0] tmp_8_fu_1331_p3;
  reg [55:0] tmp_8_reg_2838;
  wire [5:0] add_ln121_1_fu_1345_p2;
  reg [5:0] add_ln121_1_reg_2846;
  wire ap_CS_fsm_state7;
  wire [0:0] icmp_ln121_1_fu_1339_p2;
  wire [62:0] trunc_ln125_3_fu_1356_p1;
  reg [62:0] trunc_ln125_3_reg_2856;
  wire [63:0] or_ln125_1_fu_1373_p3;
  wire ap_CS_fsm_state9;
  wire [1:0] add_ln108_fu_1386_p2;
  wire ap_CS_fsm_state10;
  wire [27:0] or_ln111_2_fu_1404_p3;
  wire [0:0] icmp_ln108_fu_1380_p2;
  wire [27:0] or_ln113_2_fu_1424_p3;
  wire [55:0] tmp_16_fu_1432_p3;
  reg [55:0] tmp_16_reg_2884;
  wire [5:0] add_ln121_2_fu_1446_p2;
  reg [5:0] add_ln121_2_reg_2892;
  wire ap_CS_fsm_state11;
  wire [0:0] icmp_ln121_2_fu_1440_p2;
  wire [62:0] trunc_ln125_5_fu_1457_p1;
  reg [62:0] trunc_ln125_5_reg_2902;
  wire [63:0] or_ln125_2_fu_1474_p3;
  wire ap_CS_fsm_state13;
  wire [1:0] add_ln108_1_fu_1487_p2;
  wire ap_CS_fsm_state14;
  wire [27:0] or_ln111_3_fu_1505_p3;
  wire [0:0] icmp_ln108_1_fu_1481_p2;
  wire [27:0] or_ln113_3_fu_1525_p3;
  wire [55:0] tmp_25_fu_1533_p3;
  reg [55:0] tmp_25_reg_2930;
  wire [5:0] add_ln121_3_fu_1547_p2;
  reg [5:0] add_ln121_3_reg_2938;
  wire ap_CS_fsm_state15;
  wire [0:0] icmp_ln121_3_fu_1541_p2;
  wire [62:0] trunc_ln125_7_fu_1558_p1;
  reg [62:0] trunc_ln125_7_reg_2948;
  wire [63:0] or_ln125_3_fu_1575_p3;
  wire ap_CS_fsm_state17;
  wire [1:0] add_ln108_2_fu_1588_p2;
  wire ap_CS_fsm_state18;
  wire [27:0] or_ln111_4_fu_1606_p3;
  wire [0:0] icmp_ln108_2_fu_1582_p2;
  wire [27:0] or_ln113_4_fu_1626_p3;
  wire [55:0] tmp_28_fu_1634_p3;
  reg [55:0] tmp_28_reg_2976;
  wire [5:0] add_ln121_4_fu_1648_p2;
  reg [5:0] add_ln121_4_reg_2984;
  wire ap_CS_fsm_state19;
  wire [0:0] icmp_ln121_4_fu_1642_p2;
  wire [62:0] trunc_ln125_9_fu_1659_p1;
  reg [62:0] trunc_ln125_9_reg_2994;
  wire [63:0] or_ln125_4_fu_1676_p3;
  wire ap_CS_fsm_state21;
  wire [1:0] add_ln108_3_fu_1689_p2;
  wire ap_CS_fsm_state22;
  wire [27:0] or_ln111_5_fu_1707_p3;
  wire [0:0] icmp_ln108_3_fu_1683_p2;
  wire [27:0] or_ln113_5_fu_1727_p3;
  wire [55:0] tmp_31_fu_1735_p3;
  reg [55:0] tmp_31_reg_3022;
  wire [5:0] add_ln121_5_fu_1749_p2;
  reg [5:0] add_ln121_5_reg_3030;
  wire ap_CS_fsm_state23;
  wire [0:0] icmp_ln121_5_fu_1743_p2;
  wire [62:0] trunc_ln125_11_fu_1760_p1;
  reg [62:0] trunc_ln125_11_reg_3040;
  wire [63:0] or_ln125_5_fu_1777_p3;
  wire ap_CS_fsm_state25;
  wire [1:0] add_ln108_4_fu_1790_p2;
  wire ap_CS_fsm_state26;
  wire [27:0] or_ln111_6_fu_1808_p3;
  wire [0:0] icmp_ln108_4_fu_1784_p2;
  wire [27:0] or_ln113_6_fu_1828_p3;
  wire [55:0] tmp_34_fu_1836_p3;
  reg [55:0] tmp_34_reg_3068;
  wire [5:0] add_ln121_6_fu_1850_p2;
  reg [5:0] add_ln121_6_reg_3076;
  wire ap_CS_fsm_state27;
  wire [0:0] icmp_ln121_6_fu_1844_p2;
  wire [62:0] trunc_ln125_13_fu_1861_p1;
  reg [62:0] trunc_ln125_13_reg_3086;
  wire [63:0] or_ln125_6_fu_1878_p3;
  wire ap_CS_fsm_state29;
  wire [1:0] add_ln108_5_fu_1891_p2;
  wire ap_CS_fsm_state30;
  wire [27:0] or_ln111_7_fu_1909_p3;
  wire [0:0] icmp_ln108_5_fu_1885_p2;
  wire [27:0] or_ln113_7_fu_1929_p3;
  wire [55:0] tmp_37_fu_1937_p3;
  reg [55:0] tmp_37_reg_3114;
  wire [5:0] add_ln121_7_fu_1951_p2;
  reg [5:0] add_ln121_7_reg_3122;
  wire ap_CS_fsm_state31;
  wire [0:0] icmp_ln121_7_fu_1945_p2;
  wire [62:0] trunc_ln125_15_fu_1962_p1;
  reg [62:0] trunc_ln125_15_reg_3132;
  wire [63:0] or_ln125_7_fu_1979_p3;
  wire ap_CS_fsm_state33;
  wire [27:0] or_ln111_8_fu_1998_p3;
  wire ap_CS_fsm_state34;
  wire [0:0] ap_phi_mux_j_0_8_phi_fu_754_p4;
  wire [27:0] or_ln113_8_fu_2018_p3;
  wire [55:0] tmp_40_fu_2026_p3;
  reg [55:0] tmp_40_reg_3152;
  wire [5:0] add_ln121_8_fu_2040_p2;
  reg [5:0] add_ln121_8_reg_3160;
  wire ap_CS_fsm_state35;
  wire [0:0] icmp_ln121_8_fu_2034_p2;
  wire [62:0] trunc_ln125_17_fu_2051_p1;
  reg [62:0] trunc_ln125_17_reg_3170;
  wire [63:0] or_ln125_8_fu_2068_p3;
  wire ap_CS_fsm_state37;
  wire [1:0] add_ln108_6_fu_2081_p2;
  wire ap_CS_fsm_state38;
  wire [27:0] or_ln111_9_fu_2099_p3;
  wire [0:0] icmp_ln108_6_fu_2075_p2;
  wire [27:0] or_ln113_9_fu_2119_p3;
  wire [55:0] tmp_43_fu_2127_p3;
  reg [55:0] tmp_43_reg_3198;
  wire [5:0] add_ln121_9_fu_2141_p2;
  reg [5:0] add_ln121_9_reg_3206;
  wire ap_CS_fsm_state39;
  wire [0:0] icmp_ln121_9_fu_2135_p2;
  wire [62:0] trunc_ln125_19_fu_2152_p1;
  reg [62:0] trunc_ln125_19_reg_3216;
  wire [63:0] or_ln125_9_fu_2169_p3;
  wire ap_CS_fsm_state41;
  wire [1:0] add_ln108_7_fu_2182_p2;
  wire ap_CS_fsm_state42;
  wire [27:0] or_ln111_s_fu_2200_p3;
  wire [0:0] icmp_ln108_7_fu_2176_p2;
  wire [27:0] or_ln113_s_fu_2220_p3;
  wire [55:0] tmp_46_fu_2228_p3;
  reg [55:0] tmp_46_reg_3244;
  wire [5:0] add_ln121_10_fu_2242_p2;
  reg [5:0] add_ln121_10_reg_3252;
  wire ap_CS_fsm_state43;
  wire [0:0] icmp_ln121_10_fu_2236_p2;
  wire [62:0] trunc_ln125_21_fu_2253_p1;
  reg [62:0] trunc_ln125_21_reg_3262;
  wire [63:0] or_ln125_s_fu_2270_p3;
  wire ap_CS_fsm_state45;
  wire [1:0] add_ln108_8_fu_2283_p2;
  wire ap_CS_fsm_state46;
  wire [27:0] or_ln111_10_fu_2301_p3;
  wire [0:0] icmp_ln108_8_fu_2277_p2;
  wire [27:0] or_ln113_10_fu_2321_p3;
  wire [55:0] tmp_49_fu_2329_p3;
  reg [55:0] tmp_49_reg_3290;
  wire [5:0] add_ln121_11_fu_2343_p2;
  reg [5:0] add_ln121_11_reg_3298;
  wire ap_CS_fsm_state47;
  wire [0:0] icmp_ln121_11_fu_2337_p2;
  wire [62:0] trunc_ln125_23_fu_2354_p1;
  reg [62:0] trunc_ln125_23_reg_3308;
  wire [63:0] or_ln125_10_fu_2371_p3;
  wire ap_CS_fsm_state49;
  wire [1:0] add_ln108_9_fu_2384_p2;
  wire ap_CS_fsm_state50;
  wire [27:0] or_ln111_11_fu_2402_p3;
  wire [0:0] icmp_ln108_9_fu_2378_p2;
  wire [27:0] or_ln113_11_fu_2422_p3;
  wire [55:0] tmp_52_fu_2430_p3;
  reg [55:0] tmp_52_reg_3336;
  wire [5:0] add_ln121_12_fu_2444_p2;
  reg [5:0] add_ln121_12_reg_3344;
  wire ap_CS_fsm_state51;
  wire [0:0] icmp_ln121_12_fu_2438_p2;
  wire [62:0] trunc_ln125_25_fu_2455_p1;
  reg [62:0] trunc_ln125_25_reg_3354;
  wire [63:0] or_ln125_11_fu_2472_p3;
  wire ap_CS_fsm_state53;
  wire [1:0] add_ln108_10_fu_2485_p2;
  wire ap_CS_fsm_state54;
  wire [27:0] or_ln111_12_fu_2503_p3;
  wire [0:0] icmp_ln108_10_fu_2479_p2;
  wire [27:0] or_ln113_12_fu_2523_p3;
  wire [55:0] tmp_55_fu_2531_p3;
  reg [55:0] tmp_55_reg_3382;
  wire [5:0] add_ln121_13_fu_2545_p2;
  reg [5:0] add_ln121_13_reg_3390;
  wire ap_CS_fsm_state55;
  wire [0:0] icmp_ln121_13_fu_2539_p2;
  wire [62:0] trunc_ln125_27_fu_2556_p1;
  reg [62:0] trunc_ln125_27_reg_3400;
  wire [63:0] or_ln125_12_fu_2573_p3;
  wire ap_CS_fsm_state57;
  wire [1:0] add_ln108_11_fu_2586_p2;
  wire ap_CS_fsm_state58;
  wire [27:0] or_ln111_13_fu_2604_p3;
  wire [0:0] icmp_ln108_11_fu_2580_p2;
  wire [27:0] or_ln113_13_fu_2624_p3;
  wire [55:0] tmp_58_fu_2632_p3;
  reg [55:0] tmp_58_reg_3428;
  wire [5:0] add_ln121_14_fu_2646_p2;
  reg [5:0] add_ln121_14_reg_3436;
  wire ap_CS_fsm_state59;
  wire [0:0] icmp_ln121_14_fu_2640_p2;
  wire [62:0] trunc_ln125_29_fu_2657_p1;
  reg [62:0] trunc_ln125_29_reg_3446;
  wire [63:0] or_ln125_13_fu_2674_p3;
  wire ap_CS_fsm_state61;
  wire [27:0] or_ln111_14_fu_2693_p3;
  wire ap_CS_fsm_state62;
  wire [0:0] ap_phi_mux_j_0_15_phi_fu_1145_p4;
  wire [27:0] or_ln113_14_fu_2713_p3;
  wire [55:0] tmp_61_fu_2721_p3;
  reg [55:0] tmp_61_reg_3466;
  wire [5:0] add_ln121_15_fu_2735_p2;
  reg [5:0] add_ln121_15_reg_3474;
  wire ap_CS_fsm_state63;
  wire [0:0] icmp_ln121_15_fu_2729_p2;
  wire [62:0] trunc_ln125_31_fu_2746_p1;
  reg [62:0] trunc_ln125_31_reg_3484;
  wire [63:0] or_ln125_14_fu_2763_p3;
  wire ap_CS_fsm_state65;
  wire grp_calculationofkeys_fu_1176_ap_start;
  wire grp_calculationofkeys_fu_1176_ap_done;
  wire grp_calculationofkeys_fu_1176_ap_idle;
  wire grp_calculationofkeys_fu_1176_ap_ready;
  wire [3:0] grp_calculationofkeys_fu_1176_sub_key_address0;
  wire grp_calculationofkeys_fu_1176_sub_key_ce0;
  wire [63:0] grp_calculationofkeys_fu_1176_ap_return;
  reg [27:0] C1_reg_280;
  reg [27:0] D1_reg_290;
  reg [0:0] j_0_0_reg_300;
  reg [63:0] sub_key_load_reg_312;
  reg [5:0] j_1_0_reg_324;
  reg [27:0] C1_1_1_reg_335;
  reg [27:0] D1_1_1_reg_346;
  reg [0:0] j_0_1_reg_357;
  reg [63:0] sub_key_load_1_reg_369;
  reg [5:0] j_1_1_reg_381;
  reg [27:0] C1_1_2_reg_392;
  reg [27:0] D1_1_2_reg_403;
  reg [1:0] j_0_2_reg_414;
  reg [63:0] sub_key_load_2_reg_425;
  reg [5:0] j_1_2_reg_437;
  reg [27:0] C1_1_3_reg_448;
  reg [27:0] D1_1_3_reg_459;
  reg [1:0] j_0_3_reg_470;
  reg [63:0] sub_key_load_3_reg_481;
  reg [5:0] j_1_3_reg_493;
  reg [27:0] C1_1_4_reg_504;
  reg [27:0] D1_1_4_reg_515;
  reg [1:0] j_0_4_reg_526;
  reg [63:0] sub_key_load_4_reg_537;
  reg [5:0] j_1_4_reg_549;
  reg [27:0] C1_1_5_reg_560;
  reg [27:0] D1_1_5_reg_571;
  reg [1:0] j_0_5_reg_582;
  reg [63:0] sub_key_load_5_reg_593;
  reg [5:0] j_1_5_reg_605;
  reg [27:0] C1_1_6_reg_616;
  reg [27:0] D1_1_6_reg_627;
  reg [1:0] j_0_6_reg_638;
  reg [63:0] sub_key_load_6_reg_649;
  reg [5:0] j_1_6_reg_661;
  reg [27:0] C1_1_7_reg_672;
  reg [27:0] D1_1_7_reg_683;
  reg [1:0] j_0_7_reg_694;
  reg [63:0] sub_key_load_7_reg_705;
  reg [5:0] j_1_7_reg_717;
  reg [27:0] C1_1_8_reg_728;
  reg [27:0] D1_1_8_reg_739;
  reg [0:0] j_0_8_reg_750;
  reg [63:0] sub_key_load_8_reg_762;
  reg [5:0] j_1_8_reg_774;
  reg [27:0] C1_1_9_reg_785;
  reg [27:0] D1_1_9_reg_796;
  reg [1:0] j_0_9_reg_807;
  reg [63:0] sub_key_load_9_reg_818;
  reg [5:0] j_1_9_reg_830;
  reg [27:0] C1_1_10_reg_841;
  reg [27:0] D1_1_10_reg_852;
  reg [1:0] j_0_10_reg_863;
  reg [63:0] sub_key_load_10_reg_874;
  reg [5:0] j_1_10_reg_886;
  reg [27:0] C1_1_11_reg_897;
  reg [27:0] D1_1_11_reg_908;
  reg [1:0] j_0_11_reg_919;
  reg [63:0] sub_key_load_11_reg_930;
  reg [5:0] j_1_11_reg_942;
  reg [27:0] C1_1_12_reg_953;
  reg [27:0] D1_1_12_reg_964;
  reg [1:0] j_0_12_reg_975;
  reg [63:0] sub_key_load_12_reg_986;
  reg [5:0] j_1_12_reg_998;
  reg [27:0] C1_1_13_reg_1009;
  reg [27:0] D1_1_13_reg_1020;
  reg [1:0] j_0_13_reg_1031;
  reg [63:0] sub_key_load_13_reg_1042;
  reg [5:0] j_1_13_reg_1054;
  reg [27:0] C1_1_14_reg_1065;
  reg [27:0] D1_1_14_reg_1076;
  reg [1:0] j_0_14_reg_1087;
  reg [63:0] sub_key_load_14_reg_1098;
  reg [5:0] j_1_14_reg_1110;
  reg [27:0] C1_1_15_reg_1121;
  reg [27:0] D1_1_15_reg_1131;
  reg [0:0] j_0_15_reg_1141;
  reg [63:0] sub_key_load_15_reg_1153;
  reg [5:0] j_1_15_reg_1165;
  reg grp_calculationofkeys_fu_1176_ap_start_reg;
  wire ap_CS_fsm_state66;
  wire ap_CS_fsm_state67;
  wire [63:0] zext_ln125_fu_1262_p1;
  wire [63:0] zext_ln125_2_fu_1351_p1;
  wire [63:0] zext_ln125_4_fu_1452_p1;
  wire [63:0] zext_ln125_6_fu_1553_p1;
  wire [63:0] zext_ln125_8_fu_1654_p1;
  wire [63:0] zext_ln125_10_fu_1755_p1;
  wire [63:0] zext_ln125_12_fu_1856_p1;
  wire [63:0] zext_ln125_14_fu_1957_p1;
  wire [63:0] zext_ln125_16_fu_2046_p1;
  wire [63:0] zext_ln125_18_fu_2147_p1;
  wire [63:0] zext_ln125_20_fu_2248_p1;
  wire [63:0] zext_ln125_22_fu_2349_p1;
  wire [63:0] zext_ln125_24_fu_2450_p1;
  wire [63:0] zext_ln125_26_fu_2551_p1;
  wire [63:0] zext_ln125_28_fu_2652_p1;
  wire [63:0] zext_ln125_30_fu_2741_p1;
  wire [26:0] trunc_ln111_fu_1210_p1;
  wire [0:0] tmp_3_fu_1202_p3;
  wire [26:0] trunc_ln113_fu_1230_p1;
  wire [0:0] tmp_5_fu_1222_p3;
  wire [5:0] grp_fu_1196_p2;
  wire [55:0] zext_ln125_1_fu_1271_p1;
  wire [55:0] lshr_ln125_fu_1275_p2;
  wire [0:0] trunc_ln125_fu_1280_p1;
  wire [26:0] trunc_ln111_1_fu_1299_p1;
  wire [0:0] tmp_10_fu_1291_p3;
  wire [26:0] trunc_ln113_1_fu_1319_p1;
  wire [0:0] tmp_13_fu_1311_p3;
  wire [55:0] zext_ln125_3_fu_1360_p1;
  wire [55:0] lshr_ln125_1_fu_1364_p2;
  wire [0:0] trunc_ln125_2_fu_1369_p1;
  wire [26:0] trunc_ln111_2_fu_1400_p1;
  wire [0:0] tmp_19_fu_1392_p3;
  wire [26:0] trunc_ln113_2_fu_1420_p1;
  wire [0:0] tmp_22_fu_1412_p3;
  wire [55:0] zext_ln125_5_fu_1461_p1;
  wire [55:0] lshr_ln125_2_fu_1465_p2;
  wire [0:0] trunc_ln125_4_fu_1470_p1;
  wire [26:0] trunc_ln111_3_fu_1501_p1;
  wire [0:0] tmp_26_fu_1493_p3;
  wire [26:0] trunc_ln113_3_fu_1521_p1;
  wire [0:0] tmp_27_fu_1513_p3;
  wire [55:0] zext_ln125_7_fu_1562_p1;
  wire [55:0] lshr_ln125_3_fu_1566_p2;
  wire [0:0] trunc_ln125_6_fu_1571_p1;
  wire [26:0] trunc_ln111_4_fu_1602_p1;
  wire [0:0] tmp_29_fu_1594_p3;
  wire [26:0] trunc_ln113_4_fu_1622_p1;
  wire [0:0] tmp_30_fu_1614_p3;
  wire [55:0] zext_ln125_9_fu_1663_p1;
  wire [55:0] lshr_ln125_4_fu_1667_p2;
  wire [0:0] trunc_ln125_8_fu_1672_p1;
  wire [26:0] trunc_ln111_5_fu_1703_p1;
  wire [0:0] tmp_32_fu_1695_p3;
  wire [26:0] trunc_ln113_5_fu_1723_p1;
  wire [0:0] tmp_33_fu_1715_p3;
  wire [55:0] zext_ln125_11_fu_1764_p1;
  wire [55:0] lshr_ln125_5_fu_1768_p2;
  wire [0:0] trunc_ln125_10_fu_1773_p1;
  wire [26:0] trunc_ln111_6_fu_1804_p1;
  wire [0:0] tmp_35_fu_1796_p3;
  wire [26:0] trunc_ln113_6_fu_1824_p1;
  wire [0:0] tmp_36_fu_1816_p3;
  wire [55:0] zext_ln125_13_fu_1865_p1;
  wire [55:0] lshr_ln125_6_fu_1869_p2;
  wire [0:0] trunc_ln125_12_fu_1874_p1;
  wire [26:0] trunc_ln111_7_fu_1905_p1;
  wire [0:0] tmp_38_fu_1897_p3;
  wire [26:0] trunc_ln113_7_fu_1925_p1;
  wire [0:0] tmp_39_fu_1917_p3;
  wire [55:0] zext_ln125_15_fu_1966_p1;
  wire [55:0] lshr_ln125_7_fu_1970_p2;
  wire [0:0] trunc_ln125_14_fu_1975_p1;
  wire [26:0] trunc_ln111_8_fu_1994_p1;
  wire [0:0] tmp_41_fu_1986_p3;
  wire [26:0] trunc_ln113_8_fu_2014_p1;
  wire [0:0] tmp_42_fu_2006_p3;
  wire [55:0] zext_ln125_17_fu_2055_p1;
  wire [55:0] lshr_ln125_8_fu_2059_p2;
  wire [0:0] trunc_ln125_16_fu_2064_p1;
  wire [26:0] trunc_ln111_9_fu_2095_p1;
  wire [0:0] tmp_44_fu_2087_p3;
  wire [26:0] trunc_ln113_9_fu_2115_p1;
  wire [0:0] tmp_45_fu_2107_p3;
  wire [55:0] zext_ln125_19_fu_2156_p1;
  wire [55:0] lshr_ln125_9_fu_2160_p2;
  wire [0:0] trunc_ln125_18_fu_2165_p1;
  wire [26:0] trunc_ln111_10_fu_2196_p1;
  wire [0:0] tmp_47_fu_2188_p3;
  wire [26:0] trunc_ln113_10_fu_2216_p1;
  wire [0:0] tmp_48_fu_2208_p3;
  wire [55:0] zext_ln125_21_fu_2257_p1;
  wire [55:0] lshr_ln125_10_fu_2261_p2;
  wire [0:0] trunc_ln125_20_fu_2266_p1;
  wire [26:0] trunc_ln111_11_fu_2297_p1;
  wire [0:0] tmp_50_fu_2289_p3;
  wire [26:0] trunc_ln113_11_fu_2317_p1;
  wire [0:0] tmp_51_fu_2309_p3;
  wire [55:0] zext_ln125_23_fu_2358_p1;
  wire [55:0] lshr_ln125_11_fu_2362_p2;
  wire [0:0] trunc_ln125_22_fu_2367_p1;
  wire [26:0] trunc_ln111_12_fu_2398_p1;
  wire [0:0] tmp_53_fu_2390_p3;
  wire [26:0] trunc_ln113_12_fu_2418_p1;
  wire [0:0] tmp_54_fu_2410_p3;
  wire [55:0] zext_ln125_25_fu_2459_p1;
  wire [55:0] lshr_ln125_12_fu_2463_p2;
  wire [0:0] trunc_ln125_24_fu_2468_p1;
  wire [26:0] trunc_ln111_13_fu_2499_p1;
  wire [0:0] tmp_56_fu_2491_p3;
  wire [26:0] trunc_ln113_13_fu_2519_p1;
  wire [0:0] tmp_57_fu_2511_p3;
  wire [55:0] zext_ln125_27_fu_2560_p1;
  wire [55:0] lshr_ln125_13_fu_2564_p2;
  wire [0:0] trunc_ln125_26_fu_2569_p1;
  wire [26:0] trunc_ln111_14_fu_2600_p1;
  wire [0:0] tmp_59_fu_2592_p3;
  wire [26:0] trunc_ln113_14_fu_2620_p1;
  wire [0:0] tmp_60_fu_2612_p3;
  wire [55:0] zext_ln125_29_fu_2661_p1;
  wire [55:0] lshr_ln125_14_fu_2665_p2;
  wire [0:0] trunc_ln125_28_fu_2670_p1;
  wire [26:0] trunc_ln111_15_fu_2689_p1;
  wire [0:0] tmp_62_fu_2681_p3;
  wire [26:0] trunc_ln113_15_fu_2709_p1;
  wire [0:0] tmp_63_fu_2701_p3;
  wire [55:0] zext_ln125_31_fu_2750_p1;
  wire [55:0] lshr_ln125_15_fu_2754_p2;
  wire [0:0] trunc_ln125_30_fu_2759_p1;
  reg [63:0] ap_return_preg;
  reg [66:0] ap_NS_fsm;

  initial begin
    #0 ap_CS_fsm = 67'd1;
    #0 grp_calculationofkeys_fu_1176_ap_start_reg = 1'b0;
    #0 ap_return_preg = 64'd0;
  end


  shiftingcidi_PC2
  #(
    .DataWidth(6),
    .AddressRange(48),
    .AddressWidth(6)
  )
  PC2_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(PC2_address0),
    .ce0(PC2_ce0),
    .q0(PC2_q0)
  );


  shiftingcidi_sub_cud
  #(
    .DataWidth(64),
    .AddressRange(16),
    .AddressWidth(4)
  )
  sub_key_U
  (
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(sub_key_address0),
    .ce0(sub_key_ce0),
    .we0(sub_key_we0),
    .d0(sub_key_d0),
    .q0(sub_key_q0)
  );


  calculationofkeys
  grp_calculationofkeys_fu_1176
  (
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_calculationofkeys_fu_1176_ap_start),
    .ap_done(grp_calculationofkeys_fu_1176_ap_done),
    .ap_idle(grp_calculationofkeys_fu_1176_ap_idle),
    .ap_ready(grp_calculationofkeys_fu_1176_ap_ready),
    .L(L),
    .R(R),
    .sub_key_address0(grp_calculationofkeys_fu_1176_sub_key_address0),
    .sub_key_ce0(grp_calculationofkeys_fu_1176_sub_key_ce0),
    .sub_key_q0(sub_key_q0),
    .ap_return(grp_calculationofkeys_fu_1176_ap_return)
  );


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
      ap_CS_fsm <= ap_NS_fsm;
    end
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      ap_return_preg <= 64'd0;
    end else
      if((grp_calculationofkeys_fu_1176_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state67)) begin
        ap_return_preg <= grp_calculationofkeys_fu_1176_ap_return;
      end 
  end


  always @(posedge ap_clk) begin
    if(ap_rst == 1'b1) begin
      grp_calculationofkeys_fu_1176_ap_start_reg <= 1'b0;
    end else
      if(1'b1 == ap_CS_fsm_state66) begin
        grp_calculationofkeys_fu_1176_ap_start_reg <= 1'b1;
      end else if(grp_calculationofkeys_fu_1176_ap_ready == 1'b1) begin
        grp_calculationofkeys_fu_1176_ap_start_reg <= 1'b0;
      end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_7_fu_2176_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state42)) begin
      C1_1_10_reg_841 <= or_ln111_s_fu_2200_p3;
    end else if((icmp_ln121_9_fu_2135_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state39)) begin
      C1_1_10_reg_841 <= C1_1_9_reg_785;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_8_fu_2277_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state46)) begin
      C1_1_11_reg_897 <= or_ln111_10_fu_2301_p3;
    end else if((icmp_ln121_10_fu_2236_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state43)) begin
      C1_1_11_reg_897 <= C1_1_10_reg_841;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_9_fu_2378_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state50)) begin
      C1_1_12_reg_953 <= or_ln111_11_fu_2402_p3;
    end else if((icmp_ln121_11_fu_2337_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47)) begin
      C1_1_12_reg_953 <= C1_1_11_reg_897;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_10_fu_2479_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state54)) begin
      C1_1_13_reg_1009 <= or_ln111_12_fu_2503_p3;
    end else if((icmp_ln121_12_fu_2438_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state51)) begin
      C1_1_13_reg_1009 <= C1_1_12_reg_953;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_11_fu_2580_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state58)) begin
      C1_1_14_reg_1065 <= or_ln111_13_fu_2604_p3;
    end else if((icmp_ln121_13_fu_2539_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state55)) begin
      C1_1_14_reg_1065 <= C1_1_13_reg_1009;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state62)) begin
      C1_1_15_reg_1121 <= or_ln111_14_fu_2693_p3;
    end else if((icmp_ln121_14_fu_2640_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state59)) begin
      C1_1_15_reg_1121 <= C1_1_14_reg_1065;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      C1_1_1_reg_335 <= or_ln111_1_fu_1303_p3;
    end else if((icmp_ln121_fu_1250_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
      C1_1_1_reg_335 <= C1_reg_280;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_fu_1380_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state10)) begin
      C1_1_2_reg_392 <= or_ln111_2_fu_1404_p3;
    end else if((icmp_ln121_1_fu_1339_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
      C1_1_2_reg_392 <= C1_1_1_reg_335;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_1_fu_1481_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      C1_1_3_reg_448 <= or_ln111_3_fu_1505_p3;
    end else if((icmp_ln121_2_fu_1440_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state11)) begin
      C1_1_3_reg_448 <= C1_1_2_reg_392;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_2_fu_1582_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state18)) begin
      C1_1_4_reg_504 <= or_ln111_4_fu_1606_p3;
    end else if((icmp_ln121_3_fu_1541_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state15)) begin
      C1_1_4_reg_504 <= C1_1_3_reg_448;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_3_fu_1683_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state22)) begin
      C1_1_5_reg_560 <= or_ln111_5_fu_1707_p3;
    end else if((icmp_ln121_4_fu_1642_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state19)) begin
      C1_1_5_reg_560 <= C1_1_4_reg_504;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_4_fu_1784_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state26)) begin
      C1_1_6_reg_616 <= or_ln111_6_fu_1808_p3;
    end else if((icmp_ln121_5_fu_1743_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state23)) begin
      C1_1_6_reg_616 <= C1_1_5_reg_560;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_5_fu_1885_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state30)) begin
      C1_1_7_reg_672 <= or_ln111_7_fu_1909_p3;
    end else if((icmp_ln121_6_fu_1844_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
      C1_1_7_reg_672 <= C1_1_6_reg_616;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state34)) begin
      C1_1_8_reg_728 <= or_ln111_8_fu_1998_p3;
    end else if((icmp_ln121_7_fu_1945_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state31)) begin
      C1_1_8_reg_728 <= C1_1_7_reg_672;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_6_fu_2075_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state38)) begin
      C1_1_9_reg_785 <= or_ln111_9_fu_2099_p3;
    end else if((icmp_ln121_8_fu_2034_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state35)) begin
      C1_1_9_reg_785 <= C1_1_8_reg_728;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      C1_reg_280 <= or_ln_fu_1214_p3;
    end else if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      C1_reg_280 <= C;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_7_fu_2176_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state42)) begin
      D1_1_10_reg_852 <= or_ln113_s_fu_2220_p3;
    end else if((icmp_ln121_9_fu_2135_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state39)) begin
      D1_1_10_reg_852 <= D1_1_9_reg_796;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_8_fu_2277_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state46)) begin
      D1_1_11_reg_908 <= or_ln113_10_fu_2321_p3;
    end else if((icmp_ln121_10_fu_2236_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state43)) begin
      D1_1_11_reg_908 <= D1_1_10_reg_852;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_9_fu_2378_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state50)) begin
      D1_1_12_reg_964 <= or_ln113_11_fu_2422_p3;
    end else if((icmp_ln121_11_fu_2337_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47)) begin
      D1_1_12_reg_964 <= D1_1_11_reg_908;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_10_fu_2479_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state54)) begin
      D1_1_13_reg_1020 <= or_ln113_12_fu_2523_p3;
    end else if((icmp_ln121_12_fu_2438_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state51)) begin
      D1_1_13_reg_1020 <= D1_1_12_reg_964;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_11_fu_2580_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state58)) begin
      D1_1_14_reg_1076 <= or_ln113_13_fu_2624_p3;
    end else if((icmp_ln121_13_fu_2539_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state55)) begin
      D1_1_14_reg_1076 <= D1_1_13_reg_1020;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state62)) begin
      D1_1_15_reg_1131 <= or_ln113_14_fu_2713_p3;
    end else if((icmp_ln121_14_fu_2640_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state59)) begin
      D1_1_15_reg_1131 <= D1_1_14_reg_1076;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      D1_1_1_reg_346 <= or_ln113_1_fu_1323_p3;
    end else if((icmp_ln121_fu_1250_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
      D1_1_1_reg_346 <= D1_reg_290;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_fu_1380_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state10)) begin
      D1_1_2_reg_403 <= or_ln113_2_fu_1424_p3;
    end else if((icmp_ln121_1_fu_1339_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
      D1_1_2_reg_403 <= D1_1_1_reg_346;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_1_fu_1481_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      D1_1_3_reg_459 <= or_ln113_3_fu_1525_p3;
    end else if((icmp_ln121_2_fu_1440_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state11)) begin
      D1_1_3_reg_459 <= D1_1_2_reg_403;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_2_fu_1582_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state18)) begin
      D1_1_4_reg_515 <= or_ln113_4_fu_1626_p3;
    end else if((icmp_ln121_3_fu_1541_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state15)) begin
      D1_1_4_reg_515 <= D1_1_3_reg_459;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_3_fu_1683_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state22)) begin
      D1_1_5_reg_571 <= or_ln113_5_fu_1727_p3;
    end else if((icmp_ln121_4_fu_1642_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state19)) begin
      D1_1_5_reg_571 <= D1_1_4_reg_515;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_4_fu_1784_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state26)) begin
      D1_1_6_reg_627 <= or_ln113_6_fu_1828_p3;
    end else if((icmp_ln121_5_fu_1743_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state23)) begin
      D1_1_6_reg_627 <= D1_1_5_reg_571;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_5_fu_1885_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state30)) begin
      D1_1_7_reg_683 <= or_ln113_7_fu_1929_p3;
    end else if((icmp_ln121_6_fu_1844_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
      D1_1_7_reg_683 <= D1_1_6_reg_627;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state34)) begin
      D1_1_8_reg_739 <= or_ln113_8_fu_2018_p3;
    end else if((icmp_ln121_7_fu_1945_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state31)) begin
      D1_1_8_reg_739 <= D1_1_7_reg_683;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_6_fu_2075_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state38)) begin
      D1_1_9_reg_796 <= or_ln113_9_fu_2119_p3;
    end else if((icmp_ln121_8_fu_2034_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state35)) begin
      D1_1_9_reg_796 <= D1_1_8_reg_739;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      D1_reg_290 <= or_ln1_fu_1234_p3;
    end else if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      D1_reg_290 <= D;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state2)) begin
      j_0_0_reg_300 <= 1'd1;
    end else if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
      j_0_0_reg_300 <= 1'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_7_fu_2176_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state42)) begin
      j_0_10_reg_863 <= add_ln108_7_fu_2182_p2;
    end else if((icmp_ln121_9_fu_2135_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state39)) begin
      j_0_10_reg_863 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_8_fu_2277_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state46)) begin
      j_0_11_reg_919 <= add_ln108_8_fu_2283_p2;
    end else if((icmp_ln121_10_fu_2236_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state43)) begin
      j_0_11_reg_919 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_9_fu_2378_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state50)) begin
      j_0_12_reg_975 <= add_ln108_9_fu_2384_p2;
    end else if((icmp_ln121_11_fu_2337_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47)) begin
      j_0_12_reg_975 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_10_fu_2479_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state54)) begin
      j_0_13_reg_1031 <= add_ln108_10_fu_2485_p2;
    end else if((icmp_ln121_12_fu_2438_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state51)) begin
      j_0_13_reg_1031 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_11_fu_2580_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state58)) begin
      j_0_14_reg_1087 <= add_ln108_11_fu_2586_p2;
    end else if((icmp_ln121_13_fu_2539_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state55)) begin
      j_0_14_reg_1087 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state62)) begin
      j_0_15_reg_1141 <= 1'd1;
    end else if((icmp_ln121_14_fu_2640_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state59)) begin
      j_0_15_reg_1141 <= 1'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state6)) begin
      j_0_1_reg_357 <= 1'd1;
    end else if((icmp_ln121_fu_1250_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
      j_0_1_reg_357 <= 1'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_fu_1380_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state10)) begin
      j_0_2_reg_414 <= add_ln108_fu_1386_p2;
    end else if((icmp_ln121_1_fu_1339_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
      j_0_2_reg_414 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_1_fu_1481_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state14)) begin
      j_0_3_reg_470 <= add_ln108_1_fu_1487_p2;
    end else if((icmp_ln121_2_fu_1440_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state11)) begin
      j_0_3_reg_470 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_2_fu_1582_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state18)) begin
      j_0_4_reg_526 <= add_ln108_2_fu_1588_p2;
    end else if((icmp_ln121_3_fu_1541_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state15)) begin
      j_0_4_reg_526 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_3_fu_1683_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state22)) begin
      j_0_5_reg_582 <= add_ln108_3_fu_1689_p2;
    end else if((icmp_ln121_4_fu_1642_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state19)) begin
      j_0_5_reg_582 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_4_fu_1784_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state26)) begin
      j_0_6_reg_638 <= add_ln108_4_fu_1790_p2;
    end else if((icmp_ln121_5_fu_1743_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state23)) begin
      j_0_6_reg_638 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_5_fu_1885_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state30)) begin
      j_0_7_reg_694 <= add_ln108_5_fu_1891_p2;
    end else if((icmp_ln121_6_fu_1844_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
      j_0_7_reg_694 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd0) & (1'b1 == ap_CS_fsm_state34)) begin
      j_0_8_reg_750 <= 1'd1;
    end else if((icmp_ln121_7_fu_1945_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state31)) begin
      j_0_8_reg_750 <= 1'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_6_fu_2075_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state38)) begin
      j_0_9_reg_807 <= add_ln108_6_fu_2081_p2;
    end else if((icmp_ln121_8_fu_2034_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state35)) begin
      j_0_9_reg_807 <= 2'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      j_1_0_reg_324 <= add_ln121_reg_2808;
    end else if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      j_1_0_reg_324 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state45) begin
      j_1_10_reg_886 <= add_ln121_10_reg_3252;
    end else if((icmp_ln108_7_fu_2176_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state42)) begin
      j_1_10_reg_886 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state49) begin
      j_1_11_reg_942 <= add_ln121_11_reg_3298;
    end else if((icmp_ln108_8_fu_2277_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state46)) begin
      j_1_11_reg_942 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state53) begin
      j_1_12_reg_998 <= add_ln121_12_reg_3344;
    end else if((icmp_ln108_9_fu_2378_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state50)) begin
      j_1_12_reg_998 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state57) begin
      j_1_13_reg_1054 <= add_ln121_13_reg_3390;
    end else if((icmp_ln108_10_fu_2479_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state54)) begin
      j_1_13_reg_1054 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state61) begin
      j_1_14_reg_1110 <= add_ln121_14_reg_3436;
    end else if((icmp_ln108_11_fu_2580_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state58)) begin
      j_1_14_reg_1110 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state65) begin
      j_1_15_reg_1165 <= add_ln121_15_reg_3474;
    end else if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state62)) begin
      j_1_15_reg_1165 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      j_1_1_reg_381 <= add_ln121_1_reg_2846;
    end else if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state6)) begin
      j_1_1_reg_381 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      j_1_2_reg_437 <= add_ln121_2_reg_2892;
    end else if((icmp_ln108_fu_1380_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state10)) begin
      j_1_2_reg_437 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state17) begin
      j_1_3_reg_493 <= add_ln121_3_reg_2938;
    end else if((icmp_ln108_1_fu_1481_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
      j_1_3_reg_493 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state21) begin
      j_1_4_reg_549 <= add_ln121_4_reg_2984;
    end else if((icmp_ln108_2_fu_1582_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state18)) begin
      j_1_4_reg_549 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state25) begin
      j_1_5_reg_605 <= add_ln121_5_reg_3030;
    end else if((icmp_ln108_3_fu_1683_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state22)) begin
      j_1_5_reg_605 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state29) begin
      j_1_6_reg_661 <= add_ln121_6_reg_3076;
    end else if((icmp_ln108_4_fu_1784_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state26)) begin
      j_1_6_reg_661 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state33) begin
      j_1_7_reg_717 <= add_ln121_7_reg_3122;
    end else if((icmp_ln108_5_fu_1885_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state30)) begin
      j_1_7_reg_717 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state37) begin
      j_1_8_reg_774 <= add_ln121_8_reg_3160;
    end else if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state34)) begin
      j_1_8_reg_774 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state41) begin
      j_1_9_reg_830 <= add_ln121_9_reg_3206;
    end else if((icmp_ln108_6_fu_2075_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state38)) begin
      j_1_9_reg_830 <= 6'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state45) begin
      sub_key_load_10_reg_874 <= or_ln125_s_fu_2270_p3;
    end else if((icmp_ln108_7_fu_2176_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state42)) begin
      sub_key_load_10_reg_874 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state49) begin
      sub_key_load_11_reg_930 <= or_ln125_10_fu_2371_p3;
    end else if((icmp_ln108_8_fu_2277_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state46)) begin
      sub_key_load_11_reg_930 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state53) begin
      sub_key_load_12_reg_986 <= or_ln125_11_fu_2472_p3;
    end else if((icmp_ln108_9_fu_2378_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state50)) begin
      sub_key_load_12_reg_986 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state57) begin
      sub_key_load_13_reg_1042 <= or_ln125_12_fu_2573_p3;
    end else if((icmp_ln108_10_fu_2479_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state54)) begin
      sub_key_load_13_reg_1042 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state61) begin
      sub_key_load_14_reg_1098 <= or_ln125_13_fu_2674_p3;
    end else if((icmp_ln108_11_fu_2580_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state58)) begin
      sub_key_load_14_reg_1098 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state65) begin
      sub_key_load_15_reg_1153 <= or_ln125_14_fu_2763_p3;
    end else if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state62)) begin
      sub_key_load_15_reg_1153 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state9) begin
      sub_key_load_1_reg_369 <= or_ln125_1_fu_1373_p3;
    end else if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state6)) begin
      sub_key_load_1_reg_369 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state13) begin
      sub_key_load_2_reg_425 <= or_ln125_2_fu_1474_p3;
    end else if((icmp_ln108_fu_1380_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state10)) begin
      sub_key_load_2_reg_425 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state17) begin
      sub_key_load_3_reg_481 <= or_ln125_3_fu_1575_p3;
    end else if((icmp_ln108_1_fu_1481_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
      sub_key_load_3_reg_481 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state21) begin
      sub_key_load_4_reg_537 <= or_ln125_4_fu_1676_p3;
    end else if((icmp_ln108_2_fu_1582_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state18)) begin
      sub_key_load_4_reg_537 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state25) begin
      sub_key_load_5_reg_593 <= or_ln125_5_fu_1777_p3;
    end else if((icmp_ln108_3_fu_1683_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state22)) begin
      sub_key_load_5_reg_593 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state29) begin
      sub_key_load_6_reg_649 <= or_ln125_6_fu_1878_p3;
    end else if((icmp_ln108_4_fu_1784_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state26)) begin
      sub_key_load_6_reg_649 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state33) begin
      sub_key_load_7_reg_705 <= or_ln125_7_fu_1979_p3;
    end else if((icmp_ln108_5_fu_1885_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state30)) begin
      sub_key_load_7_reg_705 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state37) begin
      sub_key_load_8_reg_762 <= or_ln125_8_fu_2068_p3;
    end else if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state34)) begin
      sub_key_load_8_reg_762 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state41) begin
      sub_key_load_9_reg_818 <= or_ln125_9_fu_2169_p3;
    end else if((icmp_ln108_6_fu_2075_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state38)) begin
      sub_key_load_9_reg_818 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state5) begin
      sub_key_load_reg_312 <= or_ln2_fu_1284_p3;
    end else if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      sub_key_load_reg_312 <= 64'd0;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state43) begin
      add_ln121_10_reg_3252 <= add_ln121_10_fu_2242_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state47) begin
      add_ln121_11_reg_3298 <= add_ln121_11_fu_2343_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state51) begin
      add_ln121_12_reg_3344 <= add_ln121_12_fu_2444_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state55) begin
      add_ln121_13_reg_3390 <= add_ln121_13_fu_2545_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state59) begin
      add_ln121_14_reg_3436 <= add_ln121_14_fu_2646_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state63) begin
      add_ln121_15_reg_3474 <= add_ln121_15_fu_2735_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state7) begin
      add_ln121_1_reg_2846 <= add_ln121_1_fu_1345_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state11) begin
      add_ln121_2_reg_2892 <= add_ln121_2_fu_1446_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state15) begin
      add_ln121_3_reg_2938 <= add_ln121_3_fu_1547_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state19) begin
      add_ln121_4_reg_2984 <= add_ln121_4_fu_1648_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state23) begin
      add_ln121_5_reg_3030 <= add_ln121_5_fu_1749_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state27) begin
      add_ln121_6_reg_3076 <= add_ln121_6_fu_1850_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state31) begin
      add_ln121_7_reg_3122 <= add_ln121_7_fu_1951_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state35) begin
      add_ln121_8_reg_3160 <= add_ln121_8_fu_2040_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state39) begin
      add_ln121_9_reg_3206 <= add_ln121_9_fu_2141_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if(1'b1 == ap_CS_fsm_state3) begin
      add_ln121_reg_2808 <= add_ln121_fu_1256_p2;
    end 
  end


  always @(posedge ap_clk) begin
    if((1'b1 == ap_CS_fsm_state64) | (1'b1 == ap_CS_fsm_state60) | (1'b1 == ap_CS_fsm_state56) | (1'b1 == ap_CS_fsm_state52) | (1'b1 == ap_CS_fsm_state48) | (1'b1 == ap_CS_fsm_state44) | (1'b1 == ap_CS_fsm_state40) | (1'b1 == ap_CS_fsm_state36) | (1'b1 == ap_CS_fsm_state32) | (1'b1 == ap_CS_fsm_state28) | (1'b1 == ap_CS_fsm_state24) | (1'b1 == ap_CS_fsm_state20) | (1'b1 == ap_CS_fsm_state16) | (1'b1 == ap_CS_fsm_state12) | (1'b1 == ap_CS_fsm_state8) | (1'b1 == ap_CS_fsm_state4)) begin
      reg_1192 <= PC2_q0;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_fu_1380_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state10)) begin
      tmp_16_reg_2884 <= tmp_16_fu_1432_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_1_fu_1481_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
      tmp_25_reg_2930 <= tmp_25_fu_1533_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_2_fu_1582_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state18)) begin
      tmp_28_reg_2976 <= tmp_28_fu_1634_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
      tmp_2_reg_2800 <= tmp_2_fu_1242_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_3_fu_1683_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state22)) begin
      tmp_31_reg_3022 <= tmp_31_fu_1735_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_4_fu_1784_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state26)) begin
      tmp_34_reg_3068 <= tmp_34_fu_1836_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_5_fu_1885_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state30)) begin
      tmp_37_reg_3114 <= tmp_37_fu_1937_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state34)) begin
      tmp_40_reg_3152 <= tmp_40_fu_2026_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_6_fu_2075_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state38)) begin
      tmp_43_reg_3198 <= tmp_43_fu_2127_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_7_fu_2176_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state42)) begin
      tmp_46_reg_3244 <= tmp_46_fu_2228_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_8_fu_2277_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state46)) begin
      tmp_49_reg_3290 <= tmp_49_fu_2329_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_9_fu_2378_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state50)) begin
      tmp_52_reg_3336 <= tmp_52_fu_2430_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_10_fu_2479_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state54)) begin
      tmp_55_reg_3382 <= tmp_55_fu_2531_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln108_11_fu_2580_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state58)) begin
      tmp_58_reg_3428 <= tmp_58_fu_2632_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state62)) begin
      tmp_61_reg_3466 <= tmp_61_fu_2721_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state6)) begin
      tmp_8_reg_2838 <= tmp_8_fu_1331_p3;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_5_fu_1743_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state23)) begin
      trunc_ln125_11_reg_3040 <= trunc_ln125_11_fu_1760_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_6_fu_1844_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state27)) begin
      trunc_ln125_13_reg_3086 <= trunc_ln125_13_fu_1861_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_7_fu_1945_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state31)) begin
      trunc_ln125_15_reg_3132 <= trunc_ln125_15_fu_1962_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_8_fu_2034_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state35)) begin
      trunc_ln125_17_reg_3170 <= trunc_ln125_17_fu_2051_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_9_fu_2135_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state39)) begin
      trunc_ln125_19_reg_3216 <= trunc_ln125_19_fu_2152_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_fu_1250_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state3)) begin
      trunc_ln125_1_reg_2818 <= trunc_ln125_1_fu_1267_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_10_fu_2236_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state43)) begin
      trunc_ln125_21_reg_3262 <= trunc_ln125_21_fu_2253_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_11_fu_2337_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state47)) begin
      trunc_ln125_23_reg_3308 <= trunc_ln125_23_fu_2354_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_12_fu_2438_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state51)) begin
      trunc_ln125_25_reg_3354 <= trunc_ln125_25_fu_2455_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_13_fu_2539_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state55)) begin
      trunc_ln125_27_reg_3400 <= trunc_ln125_27_fu_2556_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_14_fu_2640_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state59)) begin
      trunc_ln125_29_reg_3446 <= trunc_ln125_29_fu_2657_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_15_fu_2729_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state63)) begin
      trunc_ln125_31_reg_3484 <= trunc_ln125_31_fu_2746_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_1_fu_1339_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state7)) begin
      trunc_ln125_3_reg_2856 <= trunc_ln125_3_fu_1356_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_2_fu_1440_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state11)) begin
      trunc_ln125_5_reg_2902 <= trunc_ln125_5_fu_1457_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_3_fu_1541_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state15)) begin
      trunc_ln125_7_reg_2948 <= trunc_ln125_7_fu_1558_p1;
    end 
  end


  always @(posedge ap_clk) begin
    if((icmp_ln121_4_fu_1642_p2 == 1'd0) & (1'b1 == ap_CS_fsm_state19)) begin
      trunc_ln125_9_reg_2994 <= trunc_ln125_9_fu_1659_p1;
    end 
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state63) begin
      PC2_address0 = zext_ln125_30_fu_2741_p1;
    end else if(1'b1 == ap_CS_fsm_state59) begin
      PC2_address0 = zext_ln125_28_fu_2652_p1;
    end else if(1'b1 == ap_CS_fsm_state55) begin
      PC2_address0 = zext_ln125_26_fu_2551_p1;
    end else if(1'b1 == ap_CS_fsm_state51) begin
      PC2_address0 = zext_ln125_24_fu_2450_p1;
    end else if(1'b1 == ap_CS_fsm_state47) begin
      PC2_address0 = zext_ln125_22_fu_2349_p1;
    end else if(1'b1 == ap_CS_fsm_state43) begin
      PC2_address0 = zext_ln125_20_fu_2248_p1;
    end else if(1'b1 == ap_CS_fsm_state39) begin
      PC2_address0 = zext_ln125_18_fu_2147_p1;
    end else if(1'b1 == ap_CS_fsm_state35) begin
      PC2_address0 = zext_ln125_16_fu_2046_p1;
    end else if(1'b1 == ap_CS_fsm_state31) begin
      PC2_address0 = zext_ln125_14_fu_1957_p1;
    end else if(1'b1 == ap_CS_fsm_state27) begin
      PC2_address0 = zext_ln125_12_fu_1856_p1;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      PC2_address0 = zext_ln125_10_fu_1755_p1;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      PC2_address0 = zext_ln125_8_fu_1654_p1;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      PC2_address0 = zext_ln125_6_fu_1553_p1;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      PC2_address0 = zext_ln125_4_fu_1452_p1;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      PC2_address0 = zext_ln125_2_fu_1351_p1;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      PC2_address0 = zext_ln125_fu_1262_p1;
    end else begin
      PC2_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state39) | (1'b1 == ap_CS_fsm_state35) | (1'b1 == ap_CS_fsm_state31) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state3)) begin
      PC2_ce0 = 1'b1;
    end else begin
      PC2_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1) | (grp_calculationofkeys_fu_1176_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state67)) begin
      ap_done = 1'b1;
    end else begin
      ap_done = 1'b0;
    end
  end


  always @(*) begin
    if((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)) begin
      ap_idle = 1'b1;
    end else begin
      ap_idle = 1'b0;
    end
  end


  always @(*) begin
    if((grp_calculationofkeys_fu_1176_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state67)) begin
      ap_ready = 1'b1;
    end else begin
      ap_ready = 1'b0;
    end
  end


  always @(*) begin
    if((grp_calculationofkeys_fu_1176_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state67)) begin
      ap_return = grp_calculationofkeys_fu_1176_ap_return;
    end else begin
      ap_return = ap_return_preg;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state63) begin
      sub_key_address0 = 4'd15;
    end else if(1'b1 == ap_CS_fsm_state59) begin
      sub_key_address0 = 4'd14;
    end else if(1'b1 == ap_CS_fsm_state55) begin
      sub_key_address0 = 4'd13;
    end else if(1'b1 == ap_CS_fsm_state51) begin
      sub_key_address0 = 4'd12;
    end else if(1'b1 == ap_CS_fsm_state47) begin
      sub_key_address0 = 4'd11;
    end else if(1'b1 == ap_CS_fsm_state43) begin
      sub_key_address0 = 4'd10;
    end else if(1'b1 == ap_CS_fsm_state39) begin
      sub_key_address0 = 4'd9;
    end else if(1'b1 == ap_CS_fsm_state35) begin
      sub_key_address0 = 4'd8;
    end else if(1'b1 == ap_CS_fsm_state31) begin
      sub_key_address0 = 4'd7;
    end else if(1'b1 == ap_CS_fsm_state27) begin
      sub_key_address0 = 4'd6;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      sub_key_address0 = 4'd5;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      sub_key_address0 = 4'd4;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      sub_key_address0 = 4'd3;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      sub_key_address0 = 4'd2;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      sub_key_address0 = 4'd1;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      sub_key_address0 = 4'd0;
    end else if(1'b1 == ap_CS_fsm_state67) begin
      sub_key_address0 = grp_calculationofkeys_fu_1176_sub_key_address0;
    end else begin
      sub_key_address0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state39) | (1'b1 == ap_CS_fsm_state35) | (1'b1 == ap_CS_fsm_state31) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state3)) begin
      sub_key_ce0 = 1'b1;
    end else if(1'b1 == ap_CS_fsm_state67) begin
      sub_key_ce0 = grp_calculationofkeys_fu_1176_sub_key_ce0;
    end else begin
      sub_key_ce0 = 1'b0;
    end
  end


  always @(*) begin
    if(1'b1 == ap_CS_fsm_state63) begin
      sub_key_d0 = sub_key_load_15_reg_1153;
    end else if(1'b1 == ap_CS_fsm_state59) begin
      sub_key_d0 = sub_key_load_14_reg_1098;
    end else if(1'b1 == ap_CS_fsm_state55) begin
      sub_key_d0 = sub_key_load_13_reg_1042;
    end else if(1'b1 == ap_CS_fsm_state51) begin
      sub_key_d0 = sub_key_load_12_reg_986;
    end else if(1'b1 == ap_CS_fsm_state47) begin
      sub_key_d0 = sub_key_load_11_reg_930;
    end else if(1'b1 == ap_CS_fsm_state43) begin
      sub_key_d0 = sub_key_load_10_reg_874;
    end else if(1'b1 == ap_CS_fsm_state39) begin
      sub_key_d0 = sub_key_load_9_reg_818;
    end else if(1'b1 == ap_CS_fsm_state35) begin
      sub_key_d0 = sub_key_load_8_reg_762;
    end else if(1'b1 == ap_CS_fsm_state31) begin
      sub_key_d0 = sub_key_load_7_reg_705;
    end else if(1'b1 == ap_CS_fsm_state27) begin
      sub_key_d0 = sub_key_load_6_reg_649;
    end else if(1'b1 == ap_CS_fsm_state23) begin
      sub_key_d0 = sub_key_load_5_reg_593;
    end else if(1'b1 == ap_CS_fsm_state19) begin
      sub_key_d0 = sub_key_load_4_reg_537;
    end else if(1'b1 == ap_CS_fsm_state15) begin
      sub_key_d0 = sub_key_load_3_reg_481;
    end else if(1'b1 == ap_CS_fsm_state11) begin
      sub_key_d0 = sub_key_load_2_reg_425;
    end else if(1'b1 == ap_CS_fsm_state7) begin
      sub_key_d0 = sub_key_load_1_reg_369;
    end else if(1'b1 == ap_CS_fsm_state3) begin
      sub_key_d0 = sub_key_load_reg_312;
    end else begin
      sub_key_d0 = 'bx;
    end
  end


  always @(*) begin
    if((1'b1 == ap_CS_fsm_state63) | (1'b1 == ap_CS_fsm_state59) | (1'b1 == ap_CS_fsm_state55) | (1'b1 == ap_CS_fsm_state51) | (1'b1 == ap_CS_fsm_state47) | (1'b1 == ap_CS_fsm_state43) | (1'b1 == ap_CS_fsm_state39) | (1'b1 == ap_CS_fsm_state35) | (1'b1 == ap_CS_fsm_state31) | (1'b1 == ap_CS_fsm_state27) | (1'b1 == ap_CS_fsm_state23) | (1'b1 == ap_CS_fsm_state19) | (1'b1 == ap_CS_fsm_state15) | (1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state7) | (1'b1 == ap_CS_fsm_state3)) begin
      sub_key_we0 = 1'b1;
    end else begin
      sub_key_we0 = 1'b0;
    end
  end


  always @(*) begin
    case(ap_CS_fsm)
      ap_ST_fsm_state1: begin
        if((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1)) begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end
      end
      ap_ST_fsm_state2: begin
        if((ap_phi_mux_j_0_0_phi_fu_304_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state2)) begin
          ap_NS_fsm = ap_ST_fsm_state3;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state2;
        end
      end
      ap_ST_fsm_state3: begin
        if((icmp_ln121_fu_1250_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state3)) begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state4;
        end
      end
      ap_ST_fsm_state4: begin
        ap_NS_fsm = ap_ST_fsm_state5;
      end
      ap_ST_fsm_state5: begin
        ap_NS_fsm = ap_ST_fsm_state3;
      end
      ap_ST_fsm_state6: begin
        if((ap_phi_mux_j_0_1_phi_fu_361_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state6)) begin
          ap_NS_fsm = ap_ST_fsm_state7;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state6;
        end
      end
      ap_ST_fsm_state7: begin
        if((icmp_ln121_1_fu_1339_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state7)) begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state8;
        end
      end
      ap_ST_fsm_state8: begin
        ap_NS_fsm = ap_ST_fsm_state9;
      end
      ap_ST_fsm_state9: begin
        ap_NS_fsm = ap_ST_fsm_state7;
      end
      ap_ST_fsm_state10: begin
        if((icmp_ln108_fu_1380_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state10)) begin
          ap_NS_fsm = ap_ST_fsm_state11;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state10;
        end
      end
      ap_ST_fsm_state11: begin
        if((icmp_ln121_2_fu_1440_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state11)) begin
          ap_NS_fsm = ap_ST_fsm_state14;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state12;
        end
      end
      ap_ST_fsm_state12: begin
        ap_NS_fsm = ap_ST_fsm_state13;
      end
      ap_ST_fsm_state13: begin
        ap_NS_fsm = ap_ST_fsm_state11;
      end
      ap_ST_fsm_state14: begin
        if((icmp_ln108_1_fu_1481_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state14)) begin
          ap_NS_fsm = ap_ST_fsm_state15;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state14;
        end
      end
      ap_ST_fsm_state15: begin
        if((icmp_ln121_3_fu_1541_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state15)) begin
          ap_NS_fsm = ap_ST_fsm_state18;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state16;
        end
      end
      ap_ST_fsm_state16: begin
        ap_NS_fsm = ap_ST_fsm_state17;
      end
      ap_ST_fsm_state17: begin
        ap_NS_fsm = ap_ST_fsm_state15;
      end
      ap_ST_fsm_state18: begin
        if((icmp_ln108_2_fu_1582_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state18)) begin
          ap_NS_fsm = ap_ST_fsm_state19;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state18;
        end
      end
      ap_ST_fsm_state19: begin
        if((icmp_ln121_4_fu_1642_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state19)) begin
          ap_NS_fsm = ap_ST_fsm_state22;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state20;
        end
      end
      ap_ST_fsm_state20: begin
        ap_NS_fsm = ap_ST_fsm_state21;
      end
      ap_ST_fsm_state21: begin
        ap_NS_fsm = ap_ST_fsm_state19;
      end
      ap_ST_fsm_state22: begin
        if((icmp_ln108_3_fu_1683_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state22)) begin
          ap_NS_fsm = ap_ST_fsm_state23;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state22;
        end
      end
      ap_ST_fsm_state23: begin
        if((icmp_ln121_5_fu_1743_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state23)) begin
          ap_NS_fsm = ap_ST_fsm_state26;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state24;
        end
      end
      ap_ST_fsm_state24: begin
        ap_NS_fsm = ap_ST_fsm_state25;
      end
      ap_ST_fsm_state25: begin
        ap_NS_fsm = ap_ST_fsm_state23;
      end
      ap_ST_fsm_state26: begin
        if((icmp_ln108_4_fu_1784_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state26)) begin
          ap_NS_fsm = ap_ST_fsm_state27;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state26;
        end
      end
      ap_ST_fsm_state27: begin
        if((icmp_ln121_6_fu_1844_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state27)) begin
          ap_NS_fsm = ap_ST_fsm_state30;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state28;
        end
      end
      ap_ST_fsm_state28: begin
        ap_NS_fsm = ap_ST_fsm_state29;
      end
      ap_ST_fsm_state29: begin
        ap_NS_fsm = ap_ST_fsm_state27;
      end
      ap_ST_fsm_state30: begin
        if((icmp_ln108_5_fu_1885_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state30)) begin
          ap_NS_fsm = ap_ST_fsm_state31;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state30;
        end
      end
      ap_ST_fsm_state31: begin
        if((icmp_ln121_7_fu_1945_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state31)) begin
          ap_NS_fsm = ap_ST_fsm_state34;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state32;
        end
      end
      ap_ST_fsm_state32: begin
        ap_NS_fsm = ap_ST_fsm_state33;
      end
      ap_ST_fsm_state33: begin
        ap_NS_fsm = ap_ST_fsm_state31;
      end
      ap_ST_fsm_state34: begin
        if((ap_phi_mux_j_0_8_phi_fu_754_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state34)) begin
          ap_NS_fsm = ap_ST_fsm_state35;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state34;
        end
      end
      ap_ST_fsm_state35: begin
        if((icmp_ln121_8_fu_2034_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state35)) begin
          ap_NS_fsm = ap_ST_fsm_state38;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state36;
        end
      end
      ap_ST_fsm_state36: begin
        ap_NS_fsm = ap_ST_fsm_state37;
      end
      ap_ST_fsm_state37: begin
        ap_NS_fsm = ap_ST_fsm_state35;
      end
      ap_ST_fsm_state38: begin
        if((icmp_ln108_6_fu_2075_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state38)) begin
          ap_NS_fsm = ap_ST_fsm_state39;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state38;
        end
      end
      ap_ST_fsm_state39: begin
        if((icmp_ln121_9_fu_2135_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state39)) begin
          ap_NS_fsm = ap_ST_fsm_state42;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state40;
        end
      end
      ap_ST_fsm_state40: begin
        ap_NS_fsm = ap_ST_fsm_state41;
      end
      ap_ST_fsm_state41: begin
        ap_NS_fsm = ap_ST_fsm_state39;
      end
      ap_ST_fsm_state42: begin
        if((icmp_ln108_7_fu_2176_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state42)) begin
          ap_NS_fsm = ap_ST_fsm_state43;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state42;
        end
      end
      ap_ST_fsm_state43: begin
        if((icmp_ln121_10_fu_2236_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state43)) begin
          ap_NS_fsm = ap_ST_fsm_state46;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state44;
        end
      end
      ap_ST_fsm_state44: begin
        ap_NS_fsm = ap_ST_fsm_state45;
      end
      ap_ST_fsm_state45: begin
        ap_NS_fsm = ap_ST_fsm_state43;
      end
      ap_ST_fsm_state46: begin
        if((icmp_ln108_8_fu_2277_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state46)) begin
          ap_NS_fsm = ap_ST_fsm_state47;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state46;
        end
      end
      ap_ST_fsm_state47: begin
        if((icmp_ln121_11_fu_2337_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state47)) begin
          ap_NS_fsm = ap_ST_fsm_state50;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state48;
        end
      end
      ap_ST_fsm_state48: begin
        ap_NS_fsm = ap_ST_fsm_state49;
      end
      ap_ST_fsm_state49: begin
        ap_NS_fsm = ap_ST_fsm_state47;
      end
      ap_ST_fsm_state50: begin
        if((icmp_ln108_9_fu_2378_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state50)) begin
          ap_NS_fsm = ap_ST_fsm_state51;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state50;
        end
      end
      ap_ST_fsm_state51: begin
        if((icmp_ln121_12_fu_2438_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state51)) begin
          ap_NS_fsm = ap_ST_fsm_state54;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state52;
        end
      end
      ap_ST_fsm_state52: begin
        ap_NS_fsm = ap_ST_fsm_state53;
      end
      ap_ST_fsm_state53: begin
        ap_NS_fsm = ap_ST_fsm_state51;
      end
      ap_ST_fsm_state54: begin
        if((icmp_ln108_10_fu_2479_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state54)) begin
          ap_NS_fsm = ap_ST_fsm_state55;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state54;
        end
      end
      ap_ST_fsm_state55: begin
        if((icmp_ln121_13_fu_2539_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state55)) begin
          ap_NS_fsm = ap_ST_fsm_state58;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state56;
        end
      end
      ap_ST_fsm_state56: begin
        ap_NS_fsm = ap_ST_fsm_state57;
      end
      ap_ST_fsm_state57: begin
        ap_NS_fsm = ap_ST_fsm_state55;
      end
      ap_ST_fsm_state58: begin
        if((icmp_ln108_11_fu_2580_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state58)) begin
          ap_NS_fsm = ap_ST_fsm_state59;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state58;
        end
      end
      ap_ST_fsm_state59: begin
        if((icmp_ln121_14_fu_2640_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state59)) begin
          ap_NS_fsm = ap_ST_fsm_state62;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state60;
        end
      end
      ap_ST_fsm_state60: begin
        ap_NS_fsm = ap_ST_fsm_state61;
      end
      ap_ST_fsm_state61: begin
        ap_NS_fsm = ap_ST_fsm_state59;
      end
      ap_ST_fsm_state62: begin
        if((ap_phi_mux_j_0_15_phi_fu_1145_p4 == 1'd1) & (1'b1 == ap_CS_fsm_state62)) begin
          ap_NS_fsm = ap_ST_fsm_state63;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state62;
        end
      end
      ap_ST_fsm_state63: begin
        if((icmp_ln121_15_fu_2729_p2 == 1'd1) & (1'b1 == ap_CS_fsm_state63)) begin
          ap_NS_fsm = ap_ST_fsm_state66;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state64;
        end
      end
      ap_ST_fsm_state64: begin
        ap_NS_fsm = ap_ST_fsm_state65;
      end
      ap_ST_fsm_state65: begin
        ap_NS_fsm = ap_ST_fsm_state63;
      end
      ap_ST_fsm_state66: begin
        ap_NS_fsm = ap_ST_fsm_state67;
      end
      ap_ST_fsm_state67: begin
        if((grp_calculationofkeys_fu_1176_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state67)) begin
          ap_NS_fsm = ap_ST_fsm_state1;
        end else begin
          ap_NS_fsm = ap_ST_fsm_state67;
        end
      end
      default: begin
        ap_NS_fsm = 'bx;
      end
    endcase
  end

  assign add_ln108_10_fu_2485_p2 = j_0_13_reg_1031 + 2'd1;
  assign add_ln108_11_fu_2586_p2 = j_0_14_reg_1087 + 2'd1;
  assign add_ln108_1_fu_1487_p2 = j_0_3_reg_470 + 2'd1;
  assign add_ln108_2_fu_1588_p2 = j_0_4_reg_526 + 2'd1;
  assign add_ln108_3_fu_1689_p2 = j_0_5_reg_582 + 2'd1;
  assign add_ln108_4_fu_1790_p2 = j_0_6_reg_638 + 2'd1;
  assign add_ln108_5_fu_1891_p2 = j_0_7_reg_694 + 2'd1;
  assign add_ln108_6_fu_2081_p2 = j_0_9_reg_807 + 2'd1;
  assign add_ln108_7_fu_2182_p2 = j_0_10_reg_863 + 2'd1;
  assign add_ln108_8_fu_2283_p2 = j_0_11_reg_919 + 2'd1;
  assign add_ln108_9_fu_2384_p2 = j_0_12_reg_975 + 2'd1;
  assign add_ln108_fu_1386_p2 = j_0_2_reg_414 + 2'd1;
  assign add_ln121_10_fu_2242_p2 = j_1_10_reg_886 + 6'd1;
  assign add_ln121_11_fu_2343_p2 = j_1_11_reg_942 + 6'd1;
  assign add_ln121_12_fu_2444_p2 = j_1_12_reg_998 + 6'd1;
  assign add_ln121_13_fu_2545_p2 = j_1_13_reg_1054 + 6'd1;
  assign add_ln121_14_fu_2646_p2 = j_1_14_reg_1110 + 6'd1;
  assign add_ln121_15_fu_2735_p2 = j_1_15_reg_1165 + 6'd1;
  assign add_ln121_1_fu_1345_p2 = j_1_1_reg_381 + 6'd1;
  assign add_ln121_2_fu_1446_p2 = j_1_2_reg_437 + 6'd1;
  assign add_ln121_3_fu_1547_p2 = j_1_3_reg_493 + 6'd1;
  assign add_ln121_4_fu_1648_p2 = j_1_4_reg_549 + 6'd1;
  assign add_ln121_5_fu_1749_p2 = j_1_5_reg_605 + 6'd1;
  assign add_ln121_6_fu_1850_p2 = j_1_6_reg_661 + 6'd1;
  assign add_ln121_7_fu_1951_p2 = j_1_7_reg_717 + 6'd1;
  assign add_ln121_8_fu_2040_p2 = j_1_8_reg_774 + 6'd1;
  assign add_ln121_9_fu_2141_p2 = j_1_9_reg_830 + 6'd1;
  assign add_ln121_fu_1256_p2 = j_1_0_reg_324 + 6'd1;
  assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];
  assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];
  assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];
  assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];
  assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];
  assign ap_CS_fsm_state14 = ap_CS_fsm[32'd13];
  assign ap_CS_fsm_state15 = ap_CS_fsm[32'd14];
  assign ap_CS_fsm_state16 = ap_CS_fsm[32'd15];
  assign ap_CS_fsm_state17 = ap_CS_fsm[32'd16];
  assign ap_CS_fsm_state18 = ap_CS_fsm[32'd17];
  assign ap_CS_fsm_state19 = ap_CS_fsm[32'd18];
  assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];
  assign ap_CS_fsm_state20 = ap_CS_fsm[32'd19];
  assign ap_CS_fsm_state21 = ap_CS_fsm[32'd20];
  assign ap_CS_fsm_state22 = ap_CS_fsm[32'd21];
  assign ap_CS_fsm_state23 = ap_CS_fsm[32'd22];
  assign ap_CS_fsm_state24 = ap_CS_fsm[32'd23];
  assign ap_CS_fsm_state25 = ap_CS_fsm[32'd24];
  assign ap_CS_fsm_state26 = ap_CS_fsm[32'd25];
  assign ap_CS_fsm_state27 = ap_CS_fsm[32'd26];
  assign ap_CS_fsm_state28 = ap_CS_fsm[32'd27];
  assign ap_CS_fsm_state29 = ap_CS_fsm[32'd28];
  assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];
  assign ap_CS_fsm_state30 = ap_CS_fsm[32'd29];
  assign ap_CS_fsm_state31 = ap_CS_fsm[32'd30];
  assign ap_CS_fsm_state32 = ap_CS_fsm[32'd31];
  assign ap_CS_fsm_state33 = ap_CS_fsm[32'd32];
  assign ap_CS_fsm_state34 = ap_CS_fsm[32'd33];
  assign ap_CS_fsm_state35 = ap_CS_fsm[32'd34];
  assign ap_CS_fsm_state36 = ap_CS_fsm[32'd35];
  assign ap_CS_fsm_state37 = ap_CS_fsm[32'd36];
  assign ap_CS_fsm_state38 = ap_CS_fsm[32'd37];
  assign ap_CS_fsm_state39 = ap_CS_fsm[32'd38];
  assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];
  assign ap_CS_fsm_state40 = ap_CS_fsm[32'd39];
  assign ap_CS_fsm_state41 = ap_CS_fsm[32'd40];
  assign ap_CS_fsm_state42 = ap_CS_fsm[32'd41];
  assign ap_CS_fsm_state43 = ap_CS_fsm[32'd42];
  assign ap_CS_fsm_state44 = ap_CS_fsm[32'd43];
  assign ap_CS_fsm_state45 = ap_CS_fsm[32'd44];
  assign ap_CS_fsm_state46 = ap_CS_fsm[32'd45];
  assign ap_CS_fsm_state47 = ap_CS_fsm[32'd46];
  assign ap_CS_fsm_state48 = ap_CS_fsm[32'd47];
  assign ap_CS_fsm_state49 = ap_CS_fsm[32'd48];
  assign ap_CS_fsm_state5 = ap_CS_fsm[32'd4];
  assign ap_CS_fsm_state50 = ap_CS_fsm[32'd49];
  assign ap_CS_fsm_state51 = ap_CS_fsm[32'd50];
  assign ap_CS_fsm_state52 = ap_CS_fsm[32'd51];
  assign ap_CS_fsm_state53 = ap_CS_fsm[32'd52];
  assign ap_CS_fsm_state54 = ap_CS_fsm[32'd53];
  assign ap_CS_fsm_state55 = ap_CS_fsm[32'd54];
  assign ap_CS_fsm_state56 = ap_CS_fsm[32'd55];
  assign ap_CS_fsm_state57 = ap_CS_fsm[32'd56];
  assign ap_CS_fsm_state58 = ap_CS_fsm[32'd57];
  assign ap_CS_fsm_state59 = ap_CS_fsm[32'd58];
  assign ap_CS_fsm_state6 = ap_CS_fsm[32'd5];
  assign ap_CS_fsm_state60 = ap_CS_fsm[32'd59];
  assign ap_CS_fsm_state61 = ap_CS_fsm[32'd60];
  assign ap_CS_fsm_state62 = ap_CS_fsm[32'd61];
  assign ap_CS_fsm_state63 = ap_CS_fsm[32'd62];
  assign ap_CS_fsm_state64 = ap_CS_fsm[32'd63];
  assign ap_CS_fsm_state65 = ap_CS_fsm[32'd64];
  assign ap_CS_fsm_state66 = ap_CS_fsm[32'd65];
  assign ap_CS_fsm_state67 = ap_CS_fsm[32'd66];
  assign ap_CS_fsm_state7 = ap_CS_fsm[32'd6];
  assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];
  assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];
  assign ap_phi_mux_j_0_0_phi_fu_304_p4 = j_0_0_reg_300;
  assign ap_phi_mux_j_0_15_phi_fu_1145_p4 = j_0_15_reg_1141;
  assign ap_phi_mux_j_0_1_phi_fu_361_p4 = j_0_1_reg_357;
  assign ap_phi_mux_j_0_8_phi_fu_754_p4 = j_0_8_reg_750;
  assign grp_calculationofkeys_fu_1176_ap_start = grp_calculationofkeys_fu_1176_ap_start_reg;
  assign grp_fu_1196_p2 = $signed(6'd56) - $signed(reg_1192);
  assign icmp_ln108_10_fu_2479_p2 = (j_0_13_reg_1031 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_11_fu_2580_p2 = (j_0_14_reg_1087 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_1_fu_1481_p2 = (j_0_3_reg_470 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_2_fu_1582_p2 = (j_0_4_reg_526 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_3_fu_1683_p2 = (j_0_5_reg_582 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_4_fu_1784_p2 = (j_0_6_reg_638 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_5_fu_1885_p2 = (j_0_7_reg_694 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_6_fu_2075_p2 = (j_0_9_reg_807 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_7_fu_2176_p2 = (j_0_10_reg_863 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_8_fu_2277_p2 = (j_0_11_reg_919 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_9_fu_2378_p2 = (j_0_12_reg_975 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln108_fu_1380_p2 = (j_0_2_reg_414 == 2'd2)? 1'b1 : 1'b0;
  assign icmp_ln121_10_fu_2236_p2 = (j_1_10_reg_886 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_11_fu_2337_p2 = (j_1_11_reg_942 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_12_fu_2438_p2 = (j_1_12_reg_998 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_13_fu_2539_p2 = (j_1_13_reg_1054 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_14_fu_2640_p2 = (j_1_14_reg_1110 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_15_fu_2729_p2 = (j_1_15_reg_1165 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_1_fu_1339_p2 = (j_1_1_reg_381 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_2_fu_1440_p2 = (j_1_2_reg_437 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_3_fu_1541_p2 = (j_1_3_reg_493 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_4_fu_1642_p2 = (j_1_4_reg_549 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_5_fu_1743_p2 = (j_1_5_reg_605 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_6_fu_1844_p2 = (j_1_6_reg_661 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_7_fu_1945_p2 = (j_1_7_reg_717 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_8_fu_2034_p2 = (j_1_8_reg_774 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_9_fu_2135_p2 = (j_1_9_reg_830 == 6'd48)? 1'b1 : 1'b0;
  assign icmp_ln121_fu_1250_p2 = (j_1_0_reg_324 == 6'd48)? 1'b1 : 1'b0;
  assign lshr_ln125_10_fu_2261_p2 = tmp_46_reg_3244 >> zext_ln125_21_fu_2257_p1;
  assign lshr_ln125_11_fu_2362_p2 = tmp_49_reg_3290 >> zext_ln125_23_fu_2358_p1;
  assign lshr_ln125_12_fu_2463_p2 = tmp_52_reg_3336 >> zext_ln125_25_fu_2459_p1;
  assign lshr_ln125_13_fu_2564_p2 = tmp_55_reg_3382 >> zext_ln125_27_fu_2560_p1;
  assign lshr_ln125_14_fu_2665_p2 = tmp_58_reg_3428 >> zext_ln125_29_fu_2661_p1;
  assign lshr_ln125_15_fu_2754_p2 = tmp_61_reg_3466 >> zext_ln125_31_fu_2750_p1;
  assign lshr_ln125_1_fu_1364_p2 = tmp_8_reg_2838 >> zext_ln125_3_fu_1360_p1;
  assign lshr_ln125_2_fu_1465_p2 = tmp_16_reg_2884 >> zext_ln125_5_fu_1461_p1;
  assign lshr_ln125_3_fu_1566_p2 = tmp_25_reg_2930 >> zext_ln125_7_fu_1562_p1;
  assign lshr_ln125_4_fu_1667_p2 = tmp_28_reg_2976 >> zext_ln125_9_fu_1663_p1;
  assign lshr_ln125_5_fu_1768_p2 = tmp_31_reg_3022 >> zext_ln125_11_fu_1764_p1;
  assign lshr_ln125_6_fu_1869_p2 = tmp_34_reg_3068 >> zext_ln125_13_fu_1865_p1;
  assign lshr_ln125_7_fu_1970_p2 = tmp_37_reg_3114 >> zext_ln125_15_fu_1966_p1;
  assign lshr_ln125_8_fu_2059_p2 = tmp_40_reg_3152 >> zext_ln125_17_fu_2055_p1;
  assign lshr_ln125_9_fu_2160_p2 = tmp_43_reg_3198 >> zext_ln125_19_fu_2156_p1;
  assign lshr_ln125_fu_1275_p2 = tmp_2_reg_2800 >> zext_ln125_1_fu_1271_p1;
  assign trunc_ln111_11_fu_2297_p1_temp_8 = trunc_ln111_11_fu_2297_p1 << 1'd1;
  assign trunc_ln111_11_fu_2297_p1_temp_9 = trunc_ln111_11_fu_2297_p1_temp_8 | tmp_50_fu_2289_p3;
  assign or_ln111_10_fu_2301_p3 = trunc_ln111_11_fu_2297_p1_temp_9;
  assign trunc_ln111_12_fu_2398_p1_temp_10 = trunc_ln111_12_fu_2398_p1 << 1'd1;
  assign trunc_ln111_12_fu_2398_p1_temp_11 = trunc_ln111_12_fu_2398_p1_temp_10 | tmp_53_fu_2390_p3;
  assign or_ln111_11_fu_2402_p3 = trunc_ln111_12_fu_2398_p1_temp_11;
  assign trunc_ln111_13_fu_2499_p1_temp_12 = trunc_ln111_13_fu_2499_p1 << 1'd1;
  assign trunc_ln111_13_fu_2499_p1_temp_13 = trunc_ln111_13_fu_2499_p1_temp_12 | tmp_56_fu_2491_p3;
  assign or_ln111_12_fu_2503_p3 = trunc_ln111_13_fu_2499_p1_temp_13;
  assign trunc_ln111_14_fu_2600_p1_temp_14 = trunc_ln111_14_fu_2600_p1 << 1'd1;
  assign trunc_ln111_14_fu_2600_p1_temp_15 = trunc_ln111_14_fu_2600_p1_temp_14 | tmp_59_fu_2592_p3;
  assign or_ln111_13_fu_2604_p3 = trunc_ln111_14_fu_2600_p1_temp_15;
  assign trunc_ln111_15_fu_2689_p1_temp_16 = trunc_ln111_15_fu_2689_p1 << 1'd1;
  assign trunc_ln111_15_fu_2689_p1_temp_17 = trunc_ln111_15_fu_2689_p1_temp_16 | tmp_62_fu_2681_p3;
  assign or_ln111_14_fu_2693_p3 = trunc_ln111_15_fu_2689_p1_temp_17;
  assign trunc_ln111_1_fu_1299_p1_temp_18 = trunc_ln111_1_fu_1299_p1 << 1'd1;
  assign trunc_ln111_1_fu_1299_p1_temp_19 = trunc_ln111_1_fu_1299_p1_temp_18 | tmp_10_fu_1291_p3;
  assign or_ln111_1_fu_1303_p3 = trunc_ln111_1_fu_1299_p1_temp_19;
  assign trunc_ln111_2_fu_1400_p1_temp_20 = trunc_ln111_2_fu_1400_p1 << 1'd1;
  assign trunc_ln111_2_fu_1400_p1_temp_21 = trunc_ln111_2_fu_1400_p1_temp_20 | tmp_19_fu_1392_p3;
  assign or_ln111_2_fu_1404_p3 = trunc_ln111_2_fu_1400_p1_temp_21;
  assign trunc_ln111_3_fu_1501_p1_temp_22 = trunc_ln111_3_fu_1501_p1 << 1'd1;
  assign trunc_ln111_3_fu_1501_p1_temp_23 = trunc_ln111_3_fu_1501_p1_temp_22 | tmp_26_fu_1493_p3;
  assign or_ln111_3_fu_1505_p3 = trunc_ln111_3_fu_1501_p1_temp_23;
  assign trunc_ln111_4_fu_1602_p1_temp_24 = trunc_ln111_4_fu_1602_p1 << 1'd1;
  assign trunc_ln111_4_fu_1602_p1_temp_25 = trunc_ln111_4_fu_1602_p1_temp_24 | tmp_29_fu_1594_p3;
  assign or_ln111_4_fu_1606_p3 = trunc_ln111_4_fu_1602_p1_temp_25;
  assign trunc_ln111_5_fu_1703_p1_temp_26 = trunc_ln111_5_fu_1703_p1 << 1'd1;
  assign trunc_ln111_5_fu_1703_p1_temp_27 = trunc_ln111_5_fu_1703_p1_temp_26 | tmp_32_fu_1695_p3;
  assign or_ln111_5_fu_1707_p3 = trunc_ln111_5_fu_1703_p1_temp_27;
  assign trunc_ln111_6_fu_1804_p1_temp_28 = trunc_ln111_6_fu_1804_p1 << 1'd1;
  assign trunc_ln111_6_fu_1804_p1_temp_29 = trunc_ln111_6_fu_1804_p1_temp_28 | tmp_35_fu_1796_p3;
  assign or_ln111_6_fu_1808_p3 = trunc_ln111_6_fu_1804_p1_temp_29;
  assign trunc_ln111_7_fu_1905_p1_temp_30 = trunc_ln111_7_fu_1905_p1 << 1'd1;
  assign trunc_ln111_7_fu_1905_p1_temp_31 = trunc_ln111_7_fu_1905_p1_temp_30 | tmp_38_fu_1897_p3;
  assign or_ln111_7_fu_1909_p3 = trunc_ln111_7_fu_1905_p1_temp_31;
  assign trunc_ln111_8_fu_1994_p1_temp_32 = trunc_ln111_8_fu_1994_p1 << 1'd1;
  assign trunc_ln111_8_fu_1994_p1_temp_33 = trunc_ln111_8_fu_1994_p1_temp_32 | tmp_41_fu_1986_p3;
  assign or_ln111_8_fu_1998_p3 = trunc_ln111_8_fu_1994_p1_temp_33;
  assign trunc_ln111_9_fu_2095_p1_temp_34 = trunc_ln111_9_fu_2095_p1 << 1'd1;
  assign trunc_ln111_9_fu_2095_p1_temp_35 = trunc_ln111_9_fu_2095_p1_temp_34 | tmp_44_fu_2087_p3;
  assign or_ln111_9_fu_2099_p3 = trunc_ln111_9_fu_2095_p1_temp_35;
  assign trunc_ln111_10_fu_2196_p1_temp_36 = trunc_ln111_10_fu_2196_p1 << 1'd1;
  assign trunc_ln111_10_fu_2196_p1_temp_37 = trunc_ln111_10_fu_2196_p1_temp_36 | tmp_47_fu_2188_p3;
  assign or_ln111_s_fu_2200_p3 = trunc_ln111_10_fu_2196_p1_temp_37;
  assign trunc_ln113_11_fu_2317_p1_temp_38 = trunc_ln113_11_fu_2317_p1 << 1'd1;
  assign trunc_ln113_11_fu_2317_p1_temp_39 = trunc_ln113_11_fu_2317_p1_temp_38 | tmp_51_fu_2309_p3;
  assign or_ln113_10_fu_2321_p3 = trunc_ln113_11_fu_2317_p1_temp_39;
  assign trunc_ln113_12_fu_2418_p1_temp_40 = trunc_ln113_12_fu_2418_p1 << 1'd1;
  assign trunc_ln113_12_fu_2418_p1_temp_41 = trunc_ln113_12_fu_2418_p1_temp_40 | tmp_54_fu_2410_p3;
  assign or_ln113_11_fu_2422_p3 = trunc_ln113_12_fu_2418_p1_temp_41;
  assign trunc_ln113_13_fu_2519_p1_temp_42 = trunc_ln113_13_fu_2519_p1 << 1'd1;
  assign trunc_ln113_13_fu_2519_p1_temp_43 = trunc_ln113_13_fu_2519_p1_temp_42 | tmp_57_fu_2511_p3;
  assign or_ln113_12_fu_2523_p3 = trunc_ln113_13_fu_2519_p1_temp_43;
  assign trunc_ln113_14_fu_2620_p1_temp_44 = trunc_ln113_14_fu_2620_p1 << 1'd1;
  assign trunc_ln113_14_fu_2620_p1_temp_45 = trunc_ln113_14_fu_2620_p1_temp_44 | tmp_60_fu_2612_p3;
  assign or_ln113_13_fu_2624_p3 = trunc_ln113_14_fu_2620_p1_temp_45;
  assign trunc_ln113_15_fu_2709_p1_temp_46 = trunc_ln113_15_fu_2709_p1 << 1'd1;
  assign trunc_ln113_15_fu_2709_p1_temp_47 = trunc_ln113_15_fu_2709_p1_temp_46 | tmp_63_fu_2701_p3;
  assign or_ln113_14_fu_2713_p3 = trunc_ln113_15_fu_2709_p1_temp_47;
  assign trunc_ln113_1_fu_1319_p1_temp_48 = trunc_ln113_1_fu_1319_p1 << 1'd1;
  assign trunc_ln113_1_fu_1319_p1_temp_49 = trunc_ln113_1_fu_1319_p1_temp_48 | tmp_13_fu_1311_p3;
  assign or_ln113_1_fu_1323_p3 = trunc_ln113_1_fu_1319_p1_temp_49;
  assign trunc_ln113_2_fu_1420_p1_temp_50 = trunc_ln113_2_fu_1420_p1 << 1'd1;
  assign trunc_ln113_2_fu_1420_p1_temp_51 = trunc_ln113_2_fu_1420_p1_temp_50 | tmp_22_fu_1412_p3;
  assign or_ln113_2_fu_1424_p3 = trunc_ln113_2_fu_1420_p1_temp_51;
  assign trunc_ln113_3_fu_1521_p1_temp_52 = trunc_ln113_3_fu_1521_p1 << 1'd1;
  assign trunc_ln113_3_fu_1521_p1_temp_53 = trunc_ln113_3_fu_1521_p1_temp_52 | tmp_27_fu_1513_p3;
  assign or_ln113_3_fu_1525_p3 = trunc_ln113_3_fu_1521_p1_temp_53;
  assign trunc_ln113_4_fu_1622_p1_temp_54 = trunc_ln113_4_fu_1622_p1 << 1'd1;
  assign trunc_ln113_4_fu_1622_p1_temp_55 = trunc_ln113_4_fu_1622_p1_temp_54 | tmp_30_fu_1614_p3;
  assign or_ln113_4_fu_1626_p3 = trunc_ln113_4_fu_1622_p1_temp_55;
  assign trunc_ln113_5_fu_1723_p1_temp_56 = trunc_ln113_5_fu_1723_p1 << 1'd1;
  assign trunc_ln113_5_fu_1723_p1_temp_57 = trunc_ln113_5_fu_1723_p1_temp_56 | tmp_33_fu_1715_p3;
  assign or_ln113_5_fu_1727_p3 = trunc_ln113_5_fu_1723_p1_temp_57;
  assign trunc_ln113_6_fu_1824_p1_temp_58 = trunc_ln113_6_fu_1824_p1 << 1'd1;
  assign trunc_ln113_6_fu_1824_p1_temp_59 = trunc_ln113_6_fu_1824_p1_temp_58 | tmp_36_fu_1816_p3;
  assign or_ln113_6_fu_1828_p3 = trunc_ln113_6_fu_1824_p1_temp_59;
  assign trunc_ln113_7_fu_1925_p1_temp_60 = trunc_ln113_7_fu_1925_p1 << 1'd1;
  assign trunc_ln113_7_fu_1925_p1_temp_61 = trunc_ln113_7_fu_1925_p1_temp_60 | tmp_39_fu_1917_p3;
  assign or_ln113_7_fu_1929_p3 = trunc_ln113_7_fu_1925_p1_temp_61;
  assign trunc_ln113_8_fu_2014_p1_temp_62 = trunc_ln113_8_fu_2014_p1 << 1'd1;
  assign trunc_ln113_8_fu_2014_p1_temp_63 = trunc_ln113_8_fu_2014_p1_temp_62 | tmp_42_fu_2006_p3;
  assign or_ln113_8_fu_2018_p3 = trunc_ln113_8_fu_2014_p1_temp_63;
  assign trunc_ln113_9_fu_2115_p1_temp_64 = trunc_ln113_9_fu_2115_p1 << 1'd1;
  assign trunc_ln113_9_fu_2115_p1_temp_65 = trunc_ln113_9_fu_2115_p1_temp_64 | tmp_45_fu_2107_p3;
  assign or_ln113_9_fu_2119_p3 = trunc_ln113_9_fu_2115_p1_temp_65;
  assign trunc_ln113_10_fu_2216_p1_temp_66 = trunc_ln113_10_fu_2216_p1 << 1'd1;
  assign trunc_ln113_10_fu_2216_p1_temp_67 = trunc_ln113_10_fu_2216_p1_temp_66 | tmp_48_fu_2208_p3;
  assign or_ln113_s_fu_2220_p3 = trunc_ln113_10_fu_2216_p1_temp_67;
  assign trunc_ln125_23_reg_3308_temp_68 = trunc_ln125_23_reg_3308 << 1'd1;
  assign trunc_ln125_23_reg_3308_temp_69 = trunc_ln125_23_reg_3308_temp_68 | trunc_ln125_22_fu_2367_p1;
  assign or_ln125_10_fu_2371_p3 = trunc_ln125_23_reg_3308_temp_69;
  assign trunc_ln125_25_reg_3354_temp_70 = trunc_ln125_25_reg_3354 << 1'd1;
  assign trunc_ln125_25_reg_3354_temp_71 = trunc_ln125_25_reg_3354_temp_70 | trunc_ln125_24_fu_2468_p1;
  assign or_ln125_11_fu_2472_p3 = trunc_ln125_25_reg_3354_temp_71;
  assign trunc_ln125_27_reg_3400_temp_72 = trunc_ln125_27_reg_3400 << 1'd1;
  assign trunc_ln125_27_reg_3400_temp_73 = trunc_ln125_27_reg_3400_temp_72 | trunc_ln125_26_fu_2569_p1;
  assign or_ln125_12_fu_2573_p3 = trunc_ln125_27_reg_3400_temp_73;
  assign trunc_ln125_29_reg_3446_temp_74 = trunc_ln125_29_reg_3446 << 1'd1;
  assign trunc_ln125_29_reg_3446_temp_75 = trunc_ln125_29_reg_3446_temp_74 | trunc_ln125_28_fu_2670_p1;
  assign or_ln125_13_fu_2674_p3 = trunc_ln125_29_reg_3446_temp_75;
  assign trunc_ln125_31_reg_3484_temp_76 = trunc_ln125_31_reg_3484 << 1'd1;
  assign trunc_ln125_31_reg_3484_temp_77 = trunc_ln125_31_reg_3484_temp_76 | trunc_ln125_30_fu_2759_p1;
  assign or_ln125_14_fu_2763_p3 = trunc_ln125_31_reg_3484_temp_77;
  assign trunc_ln125_3_reg_2856_temp_78 = trunc_ln125_3_reg_2856 << 1'd1;
  assign trunc_ln125_3_reg_2856_temp_79 = trunc_ln125_3_reg_2856_temp_78 | trunc_ln125_2_fu_1369_p1;
  assign or_ln125_1_fu_1373_p3 = trunc_ln125_3_reg_2856_temp_79;
  assign trunc_ln125_5_reg_2902_temp_80 = trunc_ln125_5_reg_2902 << 1'd1;
  assign trunc_ln125_5_reg_2902_temp_81 = trunc_ln125_5_reg_2902_temp_80 | trunc_ln125_4_fu_1470_p1;
  assign or_ln125_2_fu_1474_p3 = trunc_ln125_5_reg_2902_temp_81;
  assign trunc_ln125_7_reg_2948_temp_82 = trunc_ln125_7_reg_2948 << 1'd1;
  assign trunc_ln125_7_reg_2948_temp_83 = trunc_ln125_7_reg_2948_temp_82 | trunc_ln125_6_fu_1571_p1;
  assign or_ln125_3_fu_1575_p3 = trunc_ln125_7_reg_2948_temp_83;
  assign trunc_ln125_9_reg_2994_temp_84 = trunc_ln125_9_reg_2994 << 1'd1;
  assign trunc_ln125_9_reg_2994_temp_85 = trunc_ln125_9_reg_2994_temp_84 | trunc_ln125_8_fu_1672_p1;
  assign or_ln125_4_fu_1676_p3 = trunc_ln125_9_reg_2994_temp_85;
  assign trunc_ln125_11_reg_3040_temp_86 = trunc_ln125_11_reg_3040 << 1'd1;
  assign trunc_ln125_11_reg_3040_temp_87 = trunc_ln125_11_reg_3040_temp_86 | trunc_ln125_10_fu_1773_p1;
  assign or_ln125_5_fu_1777_p3 = trunc_ln125_11_reg_3040_temp_87;
  assign trunc_ln125_13_reg_3086_temp_88 = trunc_ln125_13_reg_3086 << 1'd1;
  assign trunc_ln125_13_reg_3086_temp_89 = trunc_ln125_13_reg_3086_temp_88 | trunc_ln125_12_fu_1874_p1;
  assign or_ln125_6_fu_1878_p3 = trunc_ln125_13_reg_3086_temp_89;
  assign trunc_ln125_15_reg_3132_temp_90 = trunc_ln125_15_reg_3132 << 1'd1;
  assign trunc_ln125_15_reg_3132_temp_91 = trunc_ln125_15_reg_3132_temp_90 | trunc_ln125_14_fu_1975_p1;
  assign or_ln125_7_fu_1979_p3 = trunc_ln125_15_reg_3132_temp_91;
  assign trunc_ln125_17_reg_3170_temp_92 = trunc_ln125_17_reg_3170 << 1'd1;
  assign trunc_ln125_17_reg_3170_temp_93 = trunc_ln125_17_reg_3170_temp_92 | trunc_ln125_16_fu_2064_p1;
  assign or_ln125_8_fu_2068_p3 = trunc_ln125_17_reg_3170_temp_93;
  assign trunc_ln125_19_reg_3216_temp_94 = trunc_ln125_19_reg_3216 << 1'd1;
  assign trunc_ln125_19_reg_3216_temp_95 = trunc_ln125_19_reg_3216_temp_94 | trunc_ln125_18_fu_2165_p1;
  assign or_ln125_9_fu_2169_p3 = trunc_ln125_19_reg_3216_temp_95;
  assign trunc_ln125_21_reg_3262_temp_96 = trunc_ln125_21_reg_3262 << 1'd1;
  assign trunc_ln125_21_reg_3262_temp_97 = trunc_ln125_21_reg_3262_temp_96 | trunc_ln125_20_fu_2266_p1;
  assign or_ln125_s_fu_2270_p3 = trunc_ln125_21_reg_3262_temp_97;
  assign trunc_ln113_fu_1230_p1_temp_98 = trunc_ln113_fu_1230_p1 << 1'd1;
  assign trunc_ln113_fu_1230_p1_temp_99 = trunc_ln113_fu_1230_p1_temp_98 | tmp_5_fu_1222_p3;
  assign or_ln1_fu_1234_p3 = trunc_ln113_fu_1230_p1_temp_99;
  assign trunc_ln125_1_reg_2818_temp_100 = trunc_ln125_1_reg_2818 << 1'd1;
  assign trunc_ln125_1_reg_2818_temp_101 = trunc_ln125_1_reg_2818_temp_100 | trunc_ln125_fu_1280_p1;
  assign or_ln2_fu_1284_p3 = trunc_ln125_1_reg_2818_temp_101;
  assign trunc_ln111_fu_1210_p1_temp_102 = trunc_ln111_fu_1210_p1 << 1'd1;
  assign trunc_ln111_fu_1210_p1_temp_103 = trunc_ln111_fu_1210_p1_temp_102 | tmp_3_fu_1202_p3;
  assign or_ln_fu_1214_p3 = trunc_ln111_fu_1210_p1_temp_103;
  assign C1_1_1_reg_335_temp_104 = C1_1_1_reg_335 >> 32'd27;
  assign tmp_10_fu_1291_p3 = C1_1_1_reg_335_temp_104 & 1'd1;
  assign D1_1_1_reg_346_temp_105 = D1_1_1_reg_346 >> 32'd27;
  assign tmp_13_fu_1311_p3 = D1_1_1_reg_346_temp_105 & 1'd1;
  assign C1_1_2_reg_392_temp_106 = C1_1_2_reg_392 << 1'd28;
  assign C1_1_2_reg_392_temp_107 = C1_1_2_reg_392_temp_106 | D1_1_2_reg_403;
  assign tmp_16_fu_1432_p3 = C1_1_2_reg_392_temp_107;
  assign C1_1_2_reg_392_temp_108 = C1_1_2_reg_392 >> 32'd27;
  assign tmp_19_fu_1392_p3 = C1_1_2_reg_392_temp_108 & 1'd1;
  assign D1_1_2_reg_403_temp_109 = D1_1_2_reg_403 >> 32'd27;
  assign tmp_22_fu_1412_p3 = D1_1_2_reg_403_temp_109 & 1'd1;
  assign C1_1_3_reg_448_temp_110 = C1_1_3_reg_448 << 1'd28;
  assign C1_1_3_reg_448_temp_111 = C1_1_3_reg_448_temp_110 | D1_1_3_reg_459;
  assign tmp_25_fu_1533_p3 = C1_1_3_reg_448_temp_111;
  assign C1_1_3_reg_448_temp_112 = C1_1_3_reg_448 >> 32'd27;
  assign tmp_26_fu_1493_p3 = C1_1_3_reg_448_temp_112 & 1'd1;
  assign D1_1_3_reg_459_temp_113 = D1_1_3_reg_459 >> 32'd27;
  assign tmp_27_fu_1513_p3 = D1_1_3_reg_459_temp_113 & 1'd1;
  assign C1_1_4_reg_504_temp_114 = C1_1_4_reg_504 << 1'd28;
  assign C1_1_4_reg_504_temp_115 = C1_1_4_reg_504_temp_114 | D1_1_4_reg_515;
  assign tmp_28_fu_1634_p3 = C1_1_4_reg_504_temp_115;
  assign C1_1_4_reg_504_temp_116 = C1_1_4_reg_504 >> 32'd27;
  assign tmp_29_fu_1594_p3 = C1_1_4_reg_504_temp_116 & 1'd1;
  assign C1_reg_280_temp_117 = C1_reg_280 << 1'd28;
  assign C1_reg_280_temp_118 = C1_reg_280_temp_117 | D1_reg_290;
  assign tmp_2_fu_1242_p3 = C1_reg_280_temp_118;
  assign D1_1_4_reg_515_temp_119 = D1_1_4_reg_515 >> 32'd27;
  assign tmp_30_fu_1614_p3 = D1_1_4_reg_515_temp_119 & 1'd1;
  assign C1_1_5_reg_560_temp_120 = C1_1_5_reg_560 << 1'd28;
  assign C1_1_5_reg_560_temp_121 = C1_1_5_reg_560_temp_120 | D1_1_5_reg_571;
  assign tmp_31_fu_1735_p3 = C1_1_5_reg_560_temp_121;
  assign C1_1_5_reg_560_temp_122 = C1_1_5_reg_560 >> 32'd27;
  assign tmp_32_fu_1695_p3 = C1_1_5_reg_560_temp_122 & 1'd1;
  assign D1_1_5_reg_571_temp_123 = D1_1_5_reg_571 >> 32'd27;
  assign tmp_33_fu_1715_p3 = D1_1_5_reg_571_temp_123 & 1'd1;
  assign C1_1_6_reg_616_temp_124 = C1_1_6_reg_616 << 1'd28;
  assign C1_1_6_reg_616_temp_125 = C1_1_6_reg_616_temp_124 | D1_1_6_reg_627;
  assign tmp_34_fu_1836_p3 = C1_1_6_reg_616_temp_125;
  assign C1_1_6_reg_616_temp_126 = C1_1_6_reg_616 >> 32'd27;
  assign tmp_35_fu_1796_p3 = C1_1_6_reg_616_temp_126 & 1'd1;
  assign D1_1_6_reg_627_temp_127 = D1_1_6_reg_627 >> 32'd27;
  assign tmp_36_fu_1816_p3 = D1_1_6_reg_627_temp_127 & 1'd1;
  assign C1_1_7_reg_672_temp_128 = C1_1_7_reg_672 << 1'd28;
  assign C1_1_7_reg_672_temp_129 = C1_1_7_reg_672_temp_128 | D1_1_7_reg_683;
  assign tmp_37_fu_1937_p3 = C1_1_7_reg_672_temp_129;
  assign C1_1_7_reg_672_temp_130 = C1_1_7_reg_672 >> 32'd27;
  assign tmp_38_fu_1897_p3 = C1_1_7_reg_672_temp_130 & 1'd1;
  assign D1_1_7_reg_683_temp_131 = D1_1_7_reg_683 >> 32'd27;
  assign tmp_39_fu_1917_p3 = D1_1_7_reg_683_temp_131 & 1'd1;
  assign C1_reg_280_temp_132 = C1_reg_280 >> 32'd27;
  assign tmp_3_fu_1202_p3 = C1_reg_280_temp_132 & 1'd1;
  assign C1_1_8_reg_728_temp_133 = C1_1_8_reg_728 << 1'd28;
  assign C1_1_8_reg_728_temp_134 = C1_1_8_reg_728_temp_133 | D1_1_8_reg_739;
  assign tmp_40_fu_2026_p3 = C1_1_8_reg_728_temp_134;
  assign C1_1_8_reg_728_temp_135 = C1_1_8_reg_728 >> 32'd27;
  assign tmp_41_fu_1986_p3 = C1_1_8_reg_728_temp_135 & 1'd1;
  assign D1_1_8_reg_739_temp_136 = D1_1_8_reg_739 >> 32'd27;
  assign tmp_42_fu_2006_p3 = D1_1_8_reg_739_temp_136 & 1'd1;
  assign C1_1_9_reg_785_temp_137 = C1_1_9_reg_785 << 1'd28;
  assign C1_1_9_reg_785_temp_138 = C1_1_9_reg_785_temp_137 | D1_1_9_reg_796;
  assign tmp_43_fu_2127_p3 = C1_1_9_reg_785_temp_138;
  assign C1_1_9_reg_785_temp_139 = C1_1_9_reg_785 >> 32'd27;
  assign tmp_44_fu_2087_p3 = C1_1_9_reg_785_temp_139 & 1'd1;
  assign D1_1_9_reg_796_temp_140 = D1_1_9_reg_796 >> 32'd27;
  assign tmp_45_fu_2107_p3 = D1_1_9_reg_796_temp_140 & 1'd1;
  assign C1_1_10_reg_841_temp_141 = C1_1_10_reg_841 << 1'd28;
  assign C1_1_10_reg_841_temp_142 = C1_1_10_reg_841_temp_141 | D1_1_10_reg_852;
  assign tmp_46_fu_2228_p3 = C1_1_10_reg_841_temp_142;
  assign C1_1_10_reg_841_temp_143 = C1_1_10_reg_841 >> 32'd27;
  assign tmp_47_fu_2188_p3 = C1_1_10_reg_841_temp_143 & 1'd1;
  assign D1_1_10_reg_852_temp_144 = D1_1_10_reg_852 >> 32'd27;
  assign tmp_48_fu_2208_p3 = D1_1_10_reg_852_temp_144 & 1'd1;
  assign C1_1_11_reg_897_temp_145 = C1_1_11_reg_897 << 1'd28;
  assign C1_1_11_reg_897_temp_146 = C1_1_11_reg_897_temp_145 | D1_1_11_reg_908;
  assign tmp_49_fu_2329_p3 = C1_1_11_reg_897_temp_146;
  assign C1_1_11_reg_897_temp_147 = C1_1_11_reg_897 >> 32'd27;
  assign tmp_50_fu_2289_p3 = C1_1_11_reg_897_temp_147 & 1'd1;
  assign D1_1_11_reg_908_temp_148 = D1_1_11_reg_908 >> 32'd27;
  assign tmp_51_fu_2309_p3 = D1_1_11_reg_908_temp_148 & 1'd1;
  assign C1_1_12_reg_953_temp_149 = C1_1_12_reg_953 << 1'd28;
  assign C1_1_12_reg_953_temp_150 = C1_1_12_reg_953_temp_149 | D1_1_12_reg_964;
  assign tmp_52_fu_2430_p3 = C1_1_12_reg_953_temp_150;
  assign C1_1_12_reg_953_temp_151 = C1_1_12_reg_953 >> 32'd27;
  assign tmp_53_fu_2390_p3 = C1_1_12_reg_953_temp_151 & 1'd1;
  assign D1_1_12_reg_964_temp_152 = D1_1_12_reg_964 >> 32'd27;
  assign tmp_54_fu_2410_p3 = D1_1_12_reg_964_temp_152 & 1'd1;
  assign C1_1_13_reg_1009_temp_153 = C1_1_13_reg_1009 << 1'd28;
  assign C1_1_13_reg_1009_temp_154 = C1_1_13_reg_1009_temp_153 | D1_1_13_reg_1020;
  assign tmp_55_fu_2531_p3 = C1_1_13_reg_1009_temp_154;
  assign C1_1_13_reg_1009_temp_155 = C1_1_13_reg_1009 >> 32'd27;
  assign tmp_56_fu_2491_p3 = C1_1_13_reg_1009_temp_155 & 1'd1;
  assign D1_1_13_reg_1020_temp_156 = D1_1_13_reg_1020 >> 32'd27;
  assign tmp_57_fu_2511_p3 = D1_1_13_reg_1020_temp_156 & 1'd1;
  assign C1_1_14_reg_1065_temp_157 = C1_1_14_reg_1065 << 1'd28;
  assign C1_1_14_reg_1065_temp_158 = C1_1_14_reg_1065_temp_157 | D1_1_14_reg_1076;
  assign tmp_58_fu_2632_p3 = C1_1_14_reg_1065_temp_158;
  assign C1_1_14_reg_1065_temp_159 = C1_1_14_reg_1065 >> 32'd27;
  assign tmp_59_fu_2592_p3 = C1_1_14_reg_1065_temp_159 & 1'd1;
  assign D1_reg_290_temp_160 = D1_reg_290 >> 32'd27;
  assign tmp_5_fu_1222_p3 = D1_reg_290_temp_160 & 1'd1;
  assign D1_1_14_reg_1076_temp_161 = D1_1_14_reg_1076 >> 32'd27;
  assign tmp_60_fu_2612_p3 = D1_1_14_reg_1076_temp_161 & 1'd1;
  assign C1_1_15_reg_1121_temp_162 = C1_1_15_reg_1121 << 1'd28;
  assign C1_1_15_reg_1121_temp_163 = C1_1_15_reg_1121_temp_162 | D1_1_15_reg_1131;
  assign tmp_61_fu_2721_p3 = C1_1_15_reg_1121_temp_163;
  assign C1_1_15_reg_1121_temp_164 = C1_1_15_reg_1121 >> 32'd27;
  assign tmp_62_fu_2681_p3 = C1_1_15_reg_1121_temp_164 & 1'd1;
  assign D1_1_15_reg_1131_temp_165 = D1_1_15_reg_1131 >> 32'd27;
  assign tmp_63_fu_2701_p3 = D1_1_15_reg_1131_temp_165 & 1'd1;
  assign C1_1_1_reg_335_temp_166 = C1_1_1_reg_335 << 1'd28;
  assign C1_1_1_reg_335_temp_167 = C1_1_1_reg_335_temp_166 | D1_1_1_reg_346;
  assign tmp_8_fu_1331_p3 = C1_1_1_reg_335_temp_167;
  assign trunc_ln111_10_fu_2196_p1 = (C1_1_10_reg_841 & 27'd134217727);
  assign trunc_ln111_11_fu_2297_p1 = (C1_1_11_reg_897 & 27'd134217727);
  assign trunc_ln111_12_fu_2398_p1 = (C1_1_12_reg_953 & 27'd134217727);
  assign trunc_ln111_13_fu_2499_p1 = (C1_1_13_reg_1009 & 27'd134217727);
  assign trunc_ln111_14_fu_2600_p1 = (C1_1_14_reg_1065 & 27'd134217727);
  assign trunc_ln111_15_fu_2689_p1 = (C1_1_15_reg_1121 & 27'd134217727);
  assign trunc_ln111_1_fu_1299_p1 = (C1_1_1_reg_335 & 27'd134217727);
  assign trunc_ln111_2_fu_1400_p1 = (C1_1_2_reg_392 & 27'd134217727);
  assign trunc_ln111_3_fu_1501_p1 = (C1_1_3_reg_448 & 27'd134217727);
  assign trunc_ln111_4_fu_1602_p1 = (C1_1_4_reg_504 & 27'd134217727);
  assign trunc_ln111_5_fu_1703_p1 = (C1_1_5_reg_560 & 27'd134217727);
  assign trunc_ln111_6_fu_1804_p1 = (C1_1_6_reg_616 & 27'd134217727);
  assign trunc_ln111_7_fu_1905_p1 = (C1_1_7_reg_672 & 27'd134217727);
  assign trunc_ln111_8_fu_1994_p1 = (C1_1_8_reg_728 & 27'd134217727);
  assign trunc_ln111_9_fu_2095_p1 = (C1_1_9_reg_785 & 27'd134217727);
  assign trunc_ln111_fu_1210_p1 = (C1_reg_280 & 27'd134217727);
  assign trunc_ln113_10_fu_2216_p1 = (D1_1_10_reg_852 & 27'd134217727);
  assign trunc_ln113_11_fu_2317_p1 = (D1_1_11_reg_908 & 27'd134217727);
  assign trunc_ln113_12_fu_2418_p1 = (D1_1_12_reg_964 & 27'd134217727);
  assign trunc_ln113_13_fu_2519_p1 = (D1_1_13_reg_1020 & 27'd134217727);
  assign trunc_ln113_14_fu_2620_p1 = (D1_1_14_reg_1076 & 27'd134217727);
  assign trunc_ln113_15_fu_2709_p1 = (D1_1_15_reg_1131 & 27'd134217727);
  assign trunc_ln113_1_fu_1319_p1 = (D1_1_1_reg_346 & 27'd134217727);
  assign trunc_ln113_2_fu_1420_p1 = (D1_1_2_reg_403 & 27'd134217727);
  assign trunc_ln113_3_fu_1521_p1 = (D1_1_3_reg_459 & 27'd134217727);
  assign trunc_ln113_4_fu_1622_p1 = (D1_1_4_reg_515 & 27'd134217727);
  assign trunc_ln113_5_fu_1723_p1 = (D1_1_5_reg_571 & 27'd134217727);
  assign trunc_ln113_6_fu_1824_p1 = (D1_1_6_reg_627 & 27'd134217727);
  assign trunc_ln113_7_fu_1925_p1 = (D1_1_7_reg_683 & 27'd134217727);
  assign trunc_ln113_8_fu_2014_p1 = (D1_1_8_reg_739 & 27'd134217727);
  assign trunc_ln113_9_fu_2115_p1 = (D1_1_9_reg_796 & 27'd134217727);
  assign trunc_ln113_fu_1230_p1 = (D1_reg_290 & 27'd134217727);
  assign trunc_ln125_10_fu_1773_p1 = (lshr_ln125_5_fu_1768_p2 & 1'd1);
  assign trunc_ln125_11_fu_1760_p1 = (sub_key_load_5_reg_593 & 63'd9223372036854775807);
  assign trunc_ln125_12_fu_1874_p1 = (lshr_ln125_6_fu_1869_p2 & 1'd1);
  assign trunc_ln125_13_fu_1861_p1 = (sub_key_load_6_reg_649 & 63'd9223372036854775807);
  assign trunc_ln125_14_fu_1975_p1 = (lshr_ln125_7_fu_1970_p2 & 1'd1);
  assign trunc_ln125_15_fu_1962_p1 = (sub_key_load_7_reg_705 & 63'd9223372036854775807);
  assign trunc_ln125_16_fu_2064_p1 = (lshr_ln125_8_fu_2059_p2 & 1'd1);
  assign trunc_ln125_17_fu_2051_p1 = (sub_key_load_8_reg_762 & 63'd9223372036854775807);
  assign trunc_ln125_18_fu_2165_p1 = (lshr_ln125_9_fu_2160_p2 & 1'd1);
  assign trunc_ln125_19_fu_2152_p1 = (sub_key_load_9_reg_818 & 63'd9223372036854775807);
  assign trunc_ln125_1_fu_1267_p1 = (sub_key_load_reg_312 & 63'd9223372036854775807);
  assign trunc_ln125_20_fu_2266_p1 = (lshr_ln125_10_fu_2261_p2 & 1'd1);
  assign trunc_ln125_21_fu_2253_p1 = (sub_key_load_10_reg_874 & 63'd9223372036854775807);
  assign trunc_ln125_22_fu_2367_p1 = (lshr_ln125_11_fu_2362_p2 & 1'd1);
  assign trunc_ln125_23_fu_2354_p1 = (sub_key_load_11_reg_930 & 63'd9223372036854775807);
  assign trunc_ln125_24_fu_2468_p1 = (lshr_ln125_12_fu_2463_p2 & 1'd1);
  assign trunc_ln125_25_fu_2455_p1 = (sub_key_load_12_reg_986 & 63'd9223372036854775807);
  assign trunc_ln125_26_fu_2569_p1 = (lshr_ln125_13_fu_2564_p2 & 1'd1);
  assign trunc_ln125_27_fu_2556_p1 = (sub_key_load_13_reg_1042 & 63'd9223372036854775807);
  assign trunc_ln125_28_fu_2670_p1 = (lshr_ln125_14_fu_2665_p2 & 1'd1);
  assign trunc_ln125_29_fu_2657_p1 = (sub_key_load_14_reg_1098 & 63'd9223372036854775807);
  assign trunc_ln125_2_fu_1369_p1 = (lshr_ln125_1_fu_1364_p2 & 1'd1);
  assign trunc_ln125_30_fu_2759_p1 = (lshr_ln125_15_fu_2754_p2 & 1'd1);
  assign trunc_ln125_31_fu_2746_p1 = (sub_key_load_15_reg_1153 & 63'd9223372036854775807);
  assign trunc_ln125_3_fu_1356_p1 = (sub_key_load_1_reg_369 & 63'd9223372036854775807);
  assign trunc_ln125_4_fu_1470_p1 = (lshr_ln125_2_fu_1465_p2 & 1'd1);
  assign trunc_ln125_5_fu_1457_p1 = (sub_key_load_2_reg_425 & 63'd9223372036854775807);
  assign trunc_ln125_6_fu_1571_p1 = (lshr_ln125_3_fu_1566_p2 & 1'd1);
  assign trunc_ln125_7_fu_1558_p1 = (sub_key_load_3_reg_481 & 63'd9223372036854775807);
  assign trunc_ln125_8_fu_1672_p1 = (lshr_ln125_4_fu_1667_p2 & 1'd1);
  assign trunc_ln125_9_fu_1659_p1 = (sub_key_load_4_reg_537 & 63'd9223372036854775807);
  assign trunc_ln125_fu_1280_p1 = (lshr_ln125_fu_1275_p2 & 1'd1);
  assign zext_ln125_10_fu_1755_p1 = j_1_5_reg_605;
  assign zext_ln125_11_fu_1764_p1 = grp_fu_1196_p2;
  assign zext_ln125_12_fu_1856_p1 = j_1_6_reg_661;
  assign zext_ln125_13_fu_1865_p1 = grp_fu_1196_p2;
  assign zext_ln125_14_fu_1957_p1 = j_1_7_reg_717;
  assign zext_ln125_15_fu_1966_p1 = grp_fu_1196_p2;
  assign zext_ln125_16_fu_2046_p1 = j_1_8_reg_774;
  assign zext_ln125_17_fu_2055_p1 = grp_fu_1196_p2;
  assign zext_ln125_18_fu_2147_p1 = j_1_9_reg_830;
  assign zext_ln125_19_fu_2156_p1 = grp_fu_1196_p2;
  assign zext_ln125_1_fu_1271_p1 = grp_fu_1196_p2;
  assign zext_ln125_20_fu_2248_p1 = j_1_10_reg_886;
  assign zext_ln125_21_fu_2257_p1 = grp_fu_1196_p2;
  assign zext_ln125_22_fu_2349_p1 = j_1_11_reg_942;
  assign zext_ln125_23_fu_2358_p1 = grp_fu_1196_p2;
  assign zext_ln125_24_fu_2450_p1 = j_1_12_reg_998;
  assign zext_ln125_25_fu_2459_p1 = grp_fu_1196_p2;
  assign zext_ln125_26_fu_2551_p1 = j_1_13_reg_1054;
  assign zext_ln125_27_fu_2560_p1 = grp_fu_1196_p2;
  assign zext_ln125_28_fu_2652_p1 = j_1_14_reg_1110;
  assign zext_ln125_29_fu_2661_p1 = grp_fu_1196_p2;
  assign zext_ln125_2_fu_1351_p1 = j_1_1_reg_381;
  assign zext_ln125_30_fu_2741_p1 = j_1_15_reg_1165;
  assign zext_ln125_31_fu_2750_p1 = grp_fu_1196_p2;
  assign zext_ln125_3_fu_1360_p1 = grp_fu_1196_p2;
  assign zext_ln125_4_fu_1452_p1 = j_1_2_reg_437;
  assign zext_ln125_5_fu_1461_p1 = grp_fu_1196_p2;
  assign zext_ln125_6_fu_1553_p1 = j_1_3_reg_493;
  assign zext_ln125_7_fu_1562_p1 = grp_fu_1196_p2;
  assign zext_ln125_8_fu_1654_p1 = j_1_4_reg_549;
  assign zext_ln125_9_fu_1663_p1 = grp_fu_1196_p2;
  assign zext_ln125_fu_1262_p1 = j_1_0_reg_324;

endmodule

